//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.09 Education
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18C
//Created Time: Sat Apr 22 10:08:17 2023

module Gowin_pROM_M3 (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [13:0] ad;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire [29:0] prom_inst_0_dout_w;
wire [1:0] prom_inst_0_dout;
wire [29:0] prom_inst_1_dout_w;
wire [3:2] prom_inst_1_dout;
wire [29:0] prom_inst_2_dout_w;
wire [5:4] prom_inst_2_dout;
wire [29:0] prom_inst_3_dout_w;
wire [7:6] prom_inst_3_dout;
wire [27:0] prom_inst_4_dout_w;
wire [3:0] prom_inst_4_dout;
wire [27:0] prom_inst_5_dout_w;
wire [7:4] prom_inst_5_dout;
wire [23:0] prom_inst_6_dout_w;
wire [7:0] prom_inst_6_dout;
wire dff_q_0;
wire dff_q_1;
wire mux_o_4;
wire mux_o_10;
wire mux_o_16;
wire mux_o_22;
wire mux_o_28;
wire mux_o_34;
wire mux_o_40;
wire mux_o_46;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT2 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[13])
);
defparam lut_inst_0.INIT = 4'h2;
LUT3 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[12]),
  .I2(ad[13])
);
defparam lut_inst_1.INIT = 8'h20;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ce),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13])
);
defparam lut_inst_2.INIT = 16'h2000;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[29:0],prom_inst_0_dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 2;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h134D0632252C771F0154561543363057C14BC14FC14382478A4B864F2D430C7F;
defparam prom_inst_0.INIT_RAM_01 = 256'hD5D4246E5AD1E0BBBDEE94C2FEC4C18F4F4D540F61314FD9B3BFE64953B2CEA5;
defparam prom_inst_0.INIT_RAM_02 = 256'h3724BB2B4FF343FFABDFB38EA8B136A2C4D649F6C9DD854134F4CD18671B567F;
defparam prom_inst_0.INIT_RAM_03 = 256'h13C363210E50F36A0A053B7BEE494EE5910F09341B53C6319F155F94579BD7A0;
defparam prom_inst_0.INIT_RAM_04 = 256'h07D243BBEECC0C855FFCE6DE27094DD015EA5539F02F418D3B9CD676524031C6;
defparam prom_inst_0.INIT_RAM_05 = 256'h5DC795080A58703A54EA4696DCE7B8BDE68985944EC54F898BE2CBD2080DEFBD;
defparam prom_inst_0.INIT_RAM_06 = 256'h538921548E5D286D4D517BBC088654AC5358897095D78A3CEDE5E582BA19737E;
defparam prom_inst_0.INIT_RAM_07 = 256'hBAC766255C88080670E81C9E40A1A0955353BC391B6CA022D55C563382D0F173;
defparam prom_inst_0.INIT_RAM_08 = 256'h4D9279D0A2E11055944116D488D7250D5D243924119CA0644D0464D81C640A60;
defparam prom_inst_0.INIT_RAM_09 = 256'h4C2892D0A2D144E891E8814D768464B0247E5C977075CA0A965366CB86409627;
defparam prom_inst_0.INIT_RAM_0A = 256'hD0A2F4E2289F59B96104A4251861C61451A3929E67AA0925E9D12897139D413E;
defparam prom_inst_0.INIT_RAM_0B = 256'hC20251464EA990850DA522B963C8143F91508452734579D71E7D014107A25908;
defparam prom_inst_0.INIT_RAM_0C = 256'hD85555571378DD9F054D7C8CC8FB13F90D2CEAC4710AEE14D557137B334A4686;
defparam prom_inst_0.INIT_RAM_0D = 256'hA42930239CEA3B79500152ACAB1AC6B1B57A8F8CEABA39B7E3B555696683813E;
defparam prom_inst_0.INIT_RAM_0E = 256'h954B02234837F3CDBEBFB38F5BA3EBDC953D7751951D1CC04B48C6598671CEB3;
defparam prom_inst_0.INIT_RAM_0F = 256'h6B40CF3FFBD1F6426F089D79F73FE55DBEBF9BA020004F4AEC34433910D0DBDF;
defparam prom_inst_0.INIT_RAM_10 = 256'h79D49C7C90F95515D4014B7944856117579041271C71245E54434591AB5624A4;
defparam prom_inst_0.INIT_RAM_11 = 256'h45CE42C2F1F7EFFFB456D42CC81542FFD1AC6B1AC11E695555145DB541F3FFBD;
defparam prom_inst_0.INIT_RAM_12 = 256'h8EC47BCB23441243F9E34BB0479FAA31DEF27755F742C9A0F245CC2EE57BBBC5;
defparam prom_inst_0.INIT_RAM_13 = 256'h5D865D6FFDFFFFE7547FB3B4255EEEE55DE45B65DDE75BC04596ABAFFD1729DA;
defparam prom_inst_0.INIT_RAM_14 = 256'hD6AD587EEA2F19D3B55656E65D754B529E0952F2B27235E919D155656C553557;
defparam prom_inst_0.INIT_RAM_15 = 256'hFFDB23BC92796060A8D7224B56EE45D32D76A88C24841053A967B60927992A16;
defparam prom_inst_0.INIT_RAM_16 = 256'h5D426A07C6E8AF0B8A4579D72B616291A520DFF59F95370ED7C2C33D0BCE75D4;
defparam prom_inst_0.INIT_RAM_17 = 256'h51156A4FCDD15B76631F9FCC117F17076437D92840563D950C52D05509DC12E7;
defparam prom_inst_0.INIT_RAM_18 = 256'hBCE672955CBB712055ABC77EACC1E1B6D6A70F5B516D57C48713B151290DF120;
defparam prom_inst_0.INIT_RAM_19 = 256'hADD45CE08847B8918DEF71555B47A369D3B1269555CB7519B987E3A724E04B91;
defparam prom_inst_0.INIT_RAM_1A = 256'hDA11DE05609547E7C91F907EAF957507EAF95752FA21C3957BCA550D232E4530;
defparam prom_inst_0.INIT_RAM_1B = 256'h5D6555941D6B69D7510000445D0E161445CF4B1FBB65645547F8919D047F8917;
defparam prom_inst_0.INIT_RAM_1C = 256'hEB96BA00DFA1C7B04D7EA8EF4507DAC51D67BC514C7595795D6D1E2B55D67367;
defparam prom_inst_0.INIT_RAM_1D = 256'h1572DE37BBECC36D414D7150C3837FC32DCE1818A7E56DC0AA69BAA6068AB6F4;
defparam prom_inst_0.INIT_RAM_1E = 256'h15196D4D5672841043856F556FB1D5544C55B6D29745154131D5564587455B19;
defparam prom_inst_0.INIT_RAM_1F = 256'hB08A47D046228A3BC22C5755B6D1FA081CBD607A535167AB2BFD2BED51440DB5;
defparam prom_inst_0.INIT_RAM_20 = 256'h6E7FADC54A82B8542956AB020EB194F25924424C2CBC2CBCA020202060D52930;
defparam prom_inst_0.INIT_RAM_21 = 256'hDC7DF3F0908E1B4D5C280A24EDD2C875645CFF646996D7B5A2751CBF3ACA38D8;
defparam prom_inst_0.INIT_RAM_22 = 256'h52564E78B4D4B05DAF8DCB64ECE1964E35E5915A7A1E695BD55A297106B56512;
defparam prom_inst_0.INIT_RAM_23 = 256'hF7058F17164612E03DA554B05F7D8ACE1D564D5A492D854F2473B161F65EF859;
defparam prom_inst_0.INIT_RAM_24 = 256'h2E1CA501324DB9971887106ADD6D7161F5BA5C621D5DCED86955D771A992AB74;
defparam prom_inst_0.INIT_RAM_25 = 256'h97E7546D315055558571D9411539565AC57DCD771456AD7B214CEA05C20B60E3;
defparam prom_inst_0.INIT_RAM_26 = 256'h00ADFEBD7D99005E5C57156738F4E5BF6ED595B160BF171D1FD0FE7EBECE5D55;
defparam prom_inst_0.INIT_RAM_27 = 256'h0805565C57145D9120CC31800E000801500E808C032000404A02C83620ADC000;
defparam prom_inst_0.INIT_RAM_28 = 256'hC080F9045159F5545F7156A2C56248DB5144D51558E165E71855C5467795DB6B;
defparam prom_inst_0.INIT_RAM_29 = 256'h772EC141CFDC4D5B5F741426ACB51E56535545595E4535D52514040FFA8228AE;
defparam prom_inst_0.INIT_RAM_2A = 256'hD75875717B57177D5C512551F7547D7772CC54B096B4A454A7F09742D296BFBF;
defparam prom_inst_0.INIT_RAM_2B = 256'h8C9C646436CA3E574975C49544192638543551D15751DE94F0D8AE7017CB7587;
defparam prom_inst_0.INIT_RAM_2C = 256'h416504944067261F31C76B89A99BB92BEB9B45674564625475111FDBC7F640E8;
defparam prom_inst_0.INIT_RAM_2D = 256'h59E51C7CC41C1693B1D5DAE91164224EE42648E4AE2E1C4CD6A469FDB3699B3C;
defparam prom_inst_0.INIT_RAM_2E = 256'h09C8E4E63A49B609B9DAC24D99F1CE53C5444340D0BC987C909814DD9C78701D;
defparam prom_inst_0.INIT_RAM_2F = 256'h188FBC9C34F476CF2D2FB6F521927FC1F0A9FC25AE49BC6B27E7133A405E5515;
defparam prom_inst_0.INIT_RAM_30 = 256'hA467567456745CBFC879AB847F5FA951BAD786DA77554163050360908FD188E4;
defparam prom_inst_0.INIT_RAM_31 = 256'h8C8CB0B57AACF3D04C385EF8FAEA43BFA08FFA1540E62C2E305DD3A0EDE43173;
defparam prom_inst_0.INIT_RAM_32 = 256'hA021703B69948643CADD451127E3E17B86E4135A1458242E937800004D36292C;
defparam prom_inst_0.INIT_RAM_33 = 256'h5E7E679ED91457DBD4809D023B1B042B28A2BDEC244228A249268A2970ACA010;
defparam prom_inst_0.INIT_RAM_34 = 256'hED79AFF8A07D504241B875E4A2B15F52B318AF6CA28D545451F5BC122F94DCA5;
defparam prom_inst_0.INIT_RAM_35 = 256'hEEC2BD1D55854FFBF3BEFF5319555C6715C1C70B7C6D5A64A5C550AE0AE96E4E;
defparam prom_inst_0.INIT_RAM_36 = 256'h286382F2BCC95A3B346FF19109520CFB93EEF3B902777ACE6F1B54410BF0EFF2;
defparam prom_inst_0.INIT_RAM_37 = 256'hE456D4E2428EAE3AC21B3AB38AFCEF0BDF92E793942FD5F4E15F0BC25D18E195;
defparam prom_inst_0.INIT_RAM_38 = 256'h1732C04EF260B2828EF40F3BA0EC8A6D5DD31C7A1AFE18C6EDF13A0ABEFB3B1A;
defparam prom_inst_0.INIT_RAM_39 = 256'h18A94557658675D0A17B425F5AAADF29F55D2C25459F5089F4BEE7486EEFCE44;
defparam prom_inst_0.INIT_RAM_3A = 256'h88ABDB9272FB8B62167DE6BDE49CDE2BBB6AEDED2A0D290F1D6CE5FD555D95C6;
defparam prom_inst_0.INIT_RAM_3B = 256'h557B9CA1B6890E8EA4517D38A1901529E4E14A5C44C11B023C5CEC2D4C9264E4;
defparam prom_inst_0.INIT_RAM_3C = 256'hA76074B25579ED153074B0BA9B239DF86A30A71F495C13D8974AFD85D949269E;
defparam prom_inst_0.INIT_RAM_3D = 256'h62C6C4CA5A26096786E8D30F3729F6975B29577819D5DDB742DAD0466B8F464F;
defparam prom_inst_0.INIT_RAM_3E = 256'h5394EA5F4A55DD53755931B1C28C2BB5606D17B7D773B795388ECAC0EC48A5B6;
defparam prom_inst_0.INIT_RAM_3F = 256'hBDAB31DDA46D8EFFC38CA2B28E09B8A43A8A12E2702B521F7C6EC5FCA328C2E6;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[29:0],prom_inst_1_dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 2;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h312401C28C408A0838423384A12D4098A100230C210CE5486144E1400200004C;
defparam prom_inst_1.INIT_RAM_01 = 256'h00BC080F2AD4B0D7EA47B22377A71C0568E7100BC808802550001034C10D0244;
defparam prom_inst_1.INIT_RAM_02 = 256'h913399DBCDDFA3E7874C605DE0EFF783BED30CD83F200A8D7C820E406823DE86;
defparam prom_inst_1.INIT_RAM_03 = 256'h0ACCB187CDE182FC8FC223C8F2FE0C302891189F23492D12978BDF4A2B0BE382;
defparam prom_inst_1.INIT_RAM_04 = 256'h5627C3FFFFFEF61E20024220E6844F18060E56FA262093C38CECBFBFE710922A;
defparam prom_inst_1.INIT_RAM_05 = 256'h7D1D1D3EAC73C30C7A75871C3EF997A32ECF2032CC1E660A0182A025888F040D;
defparam prom_inst_1.INIT_RAM_06 = 256'h0186196C464F108E0B47B7720A4E8042D0D0189383DA8E58EA47C76F0EA1D304;
defparam prom_inst_1.INIT_RAM_07 = 256'hFB097FB84C440D85D22D3573C3EBF0E802E22F29BFF0B2F3D583DF928CE84BBA;
defparam prom_inst_1.INIT_RAM_08 = 256'h25F5CF2184E2320460C811C8C6A18F9BAC5D0F7D7170B6F5E24C5E3D387CB7D8;
defparam prom_inst_1.INIT_RAM_09 = 256'hDD50A18942AB5E519390B0AE5F285CDE1C97EC7AB5C74C0DF4F97D7475F0D239;
defparam prom_inst_1.INIT_RAM_0A = 256'h09421B00B0A5CC5F9B2D2D6FB6FBEFBAC95BDBDEF7ACAD72F71350AB0372802D;
defparam prom_inst_1.INIT_RAM_0B = 256'hAB6B50E3AF4BD0CB83F631F22304058F7538F5D4DA0C235538DAC050C1465F0F;
defparam prom_inst_1.INIT_RAM_0C = 256'hD5135D8120FC37D7AD0344E6E7D4B01E43BA2FAA82AB3934102D90CF990BAB2B;
defparam prom_inst_1.INIT_RAM_0D = 256'hD7BE9653ACC13A8C195402E83A1E8FA1716FCFECE41B336CD3380C873CC021BA;
defparam prom_inst_1.INIT_RAM_0E = 256'hA613039B5A19C93EC6CED326CD24517500571BD2C27A7BF0991A68E368C0837C;
defparam prom_inst_1.INIT_RAM_0F = 256'h9800E7BE7BEBF96321A46EDBED3DF12EC6CCE0B13313938716D128144A5E73E5;
defparam prom_inst_1.INIT_RAM_10 = 256'h38A0989ED64C05A1520002329CE9C803B170006DC4D88D05D44404C4E99CA440;
defparam prom_inst_1.INIT_RAM_11 = 256'h11808C4E5AD96D95BF8040C4CC3D4CDF80384E23967FAA708F89EC880F7BE7BE;
defparam prom_inst_1.INIT_RAM_12 = 256'hBA49D044131009B37C2919011175219AF418139E9BE2464AD313E637333FD001;
defparam prom_inst_1.INIT_RAM_13 = 256'h046804BFD643DD70284193A6502131302808028E90240AAE70A499A1DE793C09;
defparam prom_inst_1.INIT_RAM_14 = 256'h6B2F846A0690AC0BA9DB2663231280E0AEFA01A3A3A38AE7AC0A9DB2668C9018;
defparam prom_inst_1.INIT_RAM_15 = 256'h7760B9B1CB30C02F9868137BC25102F9AFBE6B86A0BC00230C02AF0C650A6682;
defparam prom_inst_1.INIT_RAM_16 = 256'hEF4BAA018594FB4B8F1213669AF02BC4BEB2689E39279A32A1316DD72EF7BEF6;
defparam prom_inst_1.INIT_RAM_17 = 256'h35DD6A7F3BA70BE68FAD9772ACDDE20DE92A7A32201A85CCE00CF33B2C08D9BB;
defparam prom_inst_1.INIT_RAM_18 = 256'hE67313CCA27BE13F30A87B7E87BF6E02F6A1A40BE72F0224FC8F9C03DA4ABA30;
defparam prom_inst_1.INIT_RAM_19 = 256'h47731610E68C96CCC427DC4DFCCD26F33F18C1BB3044BD2CE44E8964B7D09984;
defparam prom_inst_1.INIT_RAM_1A = 256'h67A1A3813A52847BE4C7E8C0EDCC128C0EDCC1219261054C9E871334E985129B;
defparam prom_inst_1.INIT_RAM_1B = 256'hC42000ED67A93A313440002CC0E11032CF376D94943BAE9E8C5EF84028E7ED93;
defparam prom_inst_1.INIT_RAM_1C = 256'hBC9FEAE0CB6F6D013754867ABE86834008C9004486DC8EDCC72FC24BEC422BAE;
defparam prom_inst_1.INIT_RAM_1D = 256'hD55BB4891C3BCDA36064AD08EF92730764ABBDBEF53C7B51F63D8FE767DBFA62;
defparam prom_inst_1.INIT_RAM_1E = 256'h72FFE3EECBF4BD0521BDB0000D9ECAAD8FC0BC51D5A6C0FC9555B3F2D5680A48;
defparam prom_inst_1.INIT_RAM_1F = 256'h728D00F00C708A394A110AD778A7A4A47E4ED1FAC9E47C3B15162E50279EB78E;
defparam prom_inst_1.INIT_RAM_20 = 256'h490735E29FA3E1EB10D04DD246000D535E10088859621860FEF23E7276402E98;
defparam prom_inst_1.INIT_RAM_21 = 256'h0A18A130C9EBBD4C58AD8F8420C1023749EF63C9582D00B227480844098977F4;
defparam prom_inst_1.INIT_RAM_22 = 256'hC8F4903A3081BB5C2356C40105073C90B460067522FA1C96FC021AC462B65383;
defparam prom_inst_1.INIT_RAM_23 = 256'hC21D008BC010734CFCE500BB531CD6CD564016770C2CBD4C09C08007D4B0F1E2;
defparam prom_inst_1.INIT_RAM_24 = 256'hC9B0439281E600AC46BC850E640F7B09EC22B31AFE0084F664CE310400C60174;
defparam prom_inst_1.INIT_RAM_25 = 256'h0F0309EBDB5E8CC50C00B723B475543B302BF79CCBD4858CD3A00D86C12B5C1D;
defparam prom_inst_1.INIT_RAM_26 = 256'h007ACF0E3F12008434C000091BCDD0A053950DC859C0800A7170AF878D9D2F55;
defparam prom_inst_1.INIT_RAM_27 = 256'h53A9C2328C09E200212410400C002401400A801901980940AC02080F507AD000;
defparam prom_inst_1.INIT_RAM_28 = 256'hC5CA4801B6234D0236D862118E0B1A7A089E70AD630C0003CBD08D50BF6569A9;
defparam prom_inst_1.INIT_RAM_29 = 256'hAAB1804081B6270BD2BD3527A7BE85D8C9D56C06339C9EF5C270000FFE8E1A37;
defparam prom_inst_1.INIT_RAM_2A = 256'hB72159DB519D371308E78C27E089DB6141C8106327BC88418407338EA29505CD;
defparam prom_inst_1.INIT_RAM_2B = 256'hF9CEEDE1F39CA6A61B414238038C68C39E04E7A705E72E5C466576700B984211;
defparam prom_inst_1.INIT_RAM_2C = 256'h744E54E1167F7070C514435DA88BB9989A8B032110320E76546A615B599A00EB;
defparam prom_inst_1.INIT_RAM_2D = 256'hCD474F4F1455D9D3F5DD10C1657BC557157951155C7C534D34C541353446D375;
defparam prom_inst_1.INIT_RAM_2E = 256'h5EC13978407104405E1DD815D404F01CD45754BD2DF1E06C55E0F52141414FE9;
defparam prom_inst_1.INIT_RAM_2F = 256'hA711C1E16D2DADF3DD50492534C783097DC00C39101ED3F372EE147F659BB75E;
defparam prom_inst_1.INIT_RAM_30 = 256'h0021032210332FAFDC0EDCCEDDEDFCC2CCC362D100212CF15B59855D200C5137;
defparam prom_inst_1.INIT_RAM_31 = 256'hE4FC4D7D50F10CF58D437DC5D31E92262E2516B733626C293FAA9FE29ABD3C21;
defparam prom_inst_1.INIT_RAM_32 = 256'h26F896FF5DE84E6AA3C1BDA8338A2244C33842103910380C10BDC000822D3A34;
defparam prom_inst_1.INIT_RAM_33 = 256'hC2D2F8BF47A0B9F4946809C21211B72A306228A0A90C20270C70C02B04342ADC;
defparam prom_inst_1.INIT_RAM_34 = 256'h20CBFE340C3E1686A034032CCAEF4FD099080F3312A7A0B2CF2CF5DD6FC270A6;
defparam prom_inst_1.INIT_RAM_35 = 256'h388680BBC7BC841AA1A00046209D80A1909DBE3254CD780C408DACF28FBB62F6;
defparam prom_inst_1.INIT_RAM_36 = 256'h10210070381409326C81103B18B18EF4E3D30A4F464293DE3E9FCA40E02C3C09;
defparam prom_inst_1.INIT_RAM_37 = 256'hD7C5C7AF63FA3FE342F9D8DE8FA86B0300B32FE394CDCB2C012022820B3082B3;
defparam prom_inst_1.INIT_RAM_38 = 256'h108C1AA76C9003DA702EF8049CB309782A8886B48F243EFA6182B77C4B742D8F;
defparam prom_inst_1.INIT_RAM_39 = 256'h0FF8014BE32BE58FF00BFC41D9267C093763B88A4273331E4E8338C3800A86D9;
defparam prom_inst_1.INIT_RAM_3A = 256'h8CBC94E821D93F219F182FFF2FDE4A024CB93246AF231314B110E55D49EF8D2F;
defparam prom_inst_1.INIT_RAM_3B = 256'h8223E801A88DC6A24802CB10612B7508D001040B4D33207392E8C86AFCF8B4BE;
defparam prom_inst_1.INIT_RAM_3C = 256'hDE2628712AA26E85102EA3AFE0B236EE3F93F23084038946FD8F5C664FEC70C3;
defparam prom_inst_1.INIT_RAM_3D = 256'h284E47002073229F483EA2DBC309DFB44C0948CCBC8C7BA000A8E20AA9BCC246;
defparam prom_inst_1.INIT_RAM_3E = 256'h22BA2EFD4F823278E9CE32B0C2CC64C42863AC407563277F9A0D232A7684E0CF;
defparam prom_inst_1.INIT_RAM_3F = 256'hF7E92FD3ECED320011C802A384BD08EF9F08E26008FEF2BAF237BE8CA90A80B8;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[29:0],prom_inst_2_dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 2;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hE21E04024513C38C34D12749D320C004524491409140500090009000D280034B;
defparam prom_inst_2.INIT_RAM_01 = 256'h0640A4EC5D458BF0E94D45EFE36F826DF72808040FCADA8D36EE319092ABBBCA;
defparam prom_inst_2.INIT_RAM_02 = 256'hFC33F5FCD38CF575C1303C5D47E48D1392330C9624AE202AA2AA6AA4B9BEA14E;
defparam prom_inst_2.INIT_RAM_03 = 256'hBCF03644AEEB232CCFC82D8C731C8B329A831B931EDB10B1E660272DC864B0D6;
defparam prom_inst_2.INIT_RAM_04 = 256'hFAE141555555F9200AA2C7882972B0E7288284F539E238CC0EC8C32D3A9BEAA3;
defparam prom_inst_2.INIT_RAM_05 = 256'hC01033BFBCC236ACC2F0E73042B5105C22EC0C830610D01C1C079002CF70C0CE;
defparam prom_inst_2.INIT_RAM_06 = 256'h328C03130A082C78484039822C8F1CB0331A2CF1C00A2518688C8C5FCDB3342C;
defparam prom_inst_2.INIT_RAM_07 = 256'hC32F34432243CD43774C005378E8DEF34331F71C8C32363107111331C7B4C426;
defparam prom_inst_2.INIT_RAM_08 = 256'h2CD249C28798E109FB8417E3FB4F800038348D34D0D632337700374C0335B35E;
defparam prom_inst_2.INIT_RAM_09 = 256'hCC21CB8887B70021CCE1F2D8371D32C212F348B3E34DFCECD34B35BCB32CC9BF;
defparam prom_inst_2.INIT_RAM_0A = 256'h8887B24721C3488D2BACCC4FBEFBACBAE958D8C8320C8D04BB8C31C713B8412E;
defparam prom_inst_2.INIT_RAM_0B = 256'hA7E349A3A720EEC00C38FE04B9AC1857F648F0231638A2E7B8B8C001C887800F;
defparam prom_inst_2.INIT_RAM_0C = 256'h2199662C730CCCFE444C6ECF4388031C0C388F8F3BC3B8C22800432CBF43E723;
defparam prom_inst_2.INIT_RAM_0D = 256'hC83EDD31C8731E0E2556F3C0700C030218BFF5B472FF1FA0D1E0A58924E338B1;
defparam prom_inst_2.INIT_RAM_0E = 256'hE02EEB1E91BCA811E5E5C61208CE14C1CAC4E135D0C88B8D332CF0001012A321;
defparam prom_inst_2.INIT_RAM_0F = 256'h580091D75C72A0D050C401D75C6BB280E4E4D8130011308B82F2B2F0A2C73C35;
defparam prom_inst_2.INIT_RAM_10 = 256'h0E91A3E4AAECAA2A29401A0F108135300C404050E10E204107D34CCA4B10E0EC;
defparam prom_inst_2.INIT_RAM_11 = 256'h2A2FC3431E1D75D1DFE1FC33C40C835280F83E0FBC4E504430620142AE1D75C4;
defparam prom_inst_2.INIT_RAM_12 = 256'h07B1084E0C2810316CB32CC32840D03CC30FBA10B104C0FE422B6F2282ABCC2B;
defparam prom_inst_2.INIT_RAM_13 = 256'h4A114A2473E9F7328E2742E10248899288AA2A00A8AA2ADCF287321258432CA3;
defparam prom_inst_2.INIT_RAM_14 = 256'h81000E248509F8A0512184D2442821C8C7ECA1E3E3E3E248F8A312184F056251;
defparam prom_inst_2.INIT_RAM_15 = 256'hD4185210C3186083318841720A102843C830C0EA68001402CCA630DCB8E34CCA;
defparam prom_inst_2.INIT_RAM_16 = 256'h0CDFC40BE380B8635F28C87F7334B7CA039F8C3003C4E03B481025C45C7A10C8;
defparam prom_inst_2.INIT_RAM_17 = 256'h800184F00888B0207815E1717105CAEED0EAB676F0A3AFC611C78BC87CA2FFA1;
defparam prom_inst_2.INIT_RAM_18 = 256'h20F2B2CA2122232C42849E487F802C040473C0400880826C80D1FD3B243A9E70;
defparam prom_inst_2.INIT_RAM_19 = 256'hFC418328C7E2F4066CB214A00010CE04C0FC72C82B0E137F22E25F1A0F9D3349;
defparam prom_inst_2.INIT_RAM_1A = 256'h42799C068C6CE2DC806ECE25580528E2518052838CF88C063A8B28BC70DC28BC;
defparam prom_inst_2.INIT_RAM_1B = 256'h0A04C633C0532C42852000D30A12878310D1019D41CC0010E2DC244ADE6DC61A;
defparam prom_inst_2.INIT_RAM_1C = 256'hB03BE128CAC830C38CB340FA30E2770058BCC2CA2F1021006477CB1630A04F50;
defparam prom_inst_2.INIT_RAM_1D = 256'h31B4CD65E00D620886AA32EE1C379624578B0D2C358E8CE8CCB32C8B6322C962;
defparam prom_inst_2.INIT_RAM_1E = 256'h8CC00850330F02171F03C048A1FC39A5741287BDE034DB1B1BB93C2CEEC24133;
defparam prom_inst_2.INIT_RAM_1F = 256'h91E039801D35152D47FB2322C784AC89CA8137212A1A8CDDD000CF1108204C20;
defparam prom_inst_2.INIT_RAM_20 = 256'h3BECBB6C0BEFE600F5384CCF570041518CB387382EE26FE2BABEF2363670A3CA;
defparam prom_inst_2.INIT_RAM_21 = 256'h0EF88D8BC2CB2D14EBAFAF14F8A3B28C9BC8F61B1D4006547320E8EEECF123AD;
defparam prom_inst_2.INIT_RAM_22 = 256'h15C1B57F11C6C7C9B04F5C54DCD871B5D17240415C04702E309F50116658BBB4;
defparam prom_inst_2.INIT_RAM_23 = 256'hC67050F231FD800CE97CC5C73414CB013FC90C4115C9019C5BC38B1801858536;
defparam prom_inst_2.INIT_RAM_24 = 256'hCF7BD40B6FCE4E01D102D7168DD0C4E7034C064403503909C720429965CB6AE5;
defparam prom_inst_2.INIT_RAM_25 = 256'h5356230CC0813068ACEE8CBC0A21B143448C8C31E321A902B008EB20021C0F1C;
defparam prom_inst_2.INIT_RAM_26 = 256'h00C4CFE6DF93001D46CEE4A7E79C82AA08AC50D544D5CEE8C8CFA1E5E5C88C6C;
defparam prom_inst_2.INIT_RAM_27 = 256'h4FB110C1312228200229242000001400E00D0012013809901381DC0380C4C000;
defparam prom_inst_2.INIT_RAM_28 = 256'h3D8000058780134C000ECD0000D32C0B4C2004004064A8A9E034005B33F13353;
defparam prom_inst_2.INIT_RAM_29 = 256'hEA220186000380400A31C9CD3F326120202C4D30CB2200C93480000FFE9EAC2E;
defparam prom_inst_2.INIT_RAM_2A = 256'h0483F1007F1044844008210C14020048803B2822C320A7A9CAA7280B92A56CE1;
defparam prom_inst_2.INIT_RAM_2B = 256'hCEDCDCDFE3C8F404946A188500CCB0DB10840C88840801262D1A17300054581C;
defparam prom_inst_2.INIT_RAM_2C = 256'h00101501050001010451140099A988B82133322222111A76447046BA933000EA;
defparam prom_inst_2.INIT_RAM_2D = 256'h0010001015400004050145144000000040400540014144114115114045101441;
defparam prom_inst_2.INIT_RAM_2E = 256'h5015420155045554405018140440010014100501410105010105015445151000;
defparam prom_inst_2.INIT_RAM_2F = 256'h4000110202420000001141004404141400155140441007F401AA454006400080;
defparam prom_inst_2.INIT_RAM_30 = 256'h32111000003336B67A2444477464575B646A894B130336628090190240406540;
defparam prom_inst_2.INIT_RAM_31 = 256'h7878700055015104381041000440E4C0408044C88CCCCC047FF4B9788AA6AB1A;
defparam prom_inst_2.INIT_RAM_32 = 256'hA916E37E4EC00EB603486242018AFAA203BC22AC0404AA3BC8BC0C0004121030;
defparam prom_inst_2.INIT_RAM_33 = 256'h6212348F484AC79CB288EBCE3A38BB2A28A1CC50A70A28A904504A19069CF2EC;
defparam prom_inst_2.INIT_RAM_34 = 256'hD208FA3CAB5F5F4AD2E34822CED85222BB2CAFA411E86AC30800C8ECC7DA88A9;
defparam prom_inst_2.INIT_RAM_35 = 256'hBA8A70C50C71EDB562ABBA9E3A5208E69DA4622AF4785530AD4102FBAF94DCF5;
defparam prom_inst_2.INIT_RAM_36 = 256'h18E38EA3ED8C241A20EBB2DC28025CEAE9ABA2EC0AA6510F409412419EEEBAA3;
defparam prom_inst_2.INIT_RAM_37 = 256'hC1C1155F3FD4FF53CF7372C52FA8A83E208B23C1887AA800E3BA2A8A0C38E394;
defparam prom_inst_2.INIT_RAM_38 = 256'h0B51AB2F1053C8CB45A50AD2F2F82F7938B16AD8EFA48F1FD6BB3B13E8D8FCEF;
defparam prom_inst_2.INIT_RAM_39 = 256'h8CF501230C912980F0631BBB334CB22A909808AC25C981ED472BB1C7155A8A00;
defparam prom_inst_2.INIT_RAM_3A = 256'h2DFE8206A00A7D91155923C823D2C72A6673B94EBF2E298C4C086821210C32B0;
defparam prom_inst_2.INIT_RAM_3B = 256'h2C1EC8A3A627CE5107BB0038A38BBE28F8E38ACCC7331C0B3108E8A8FFDD3337;
defparam prom_inst_2.INIT_RAM_3C = 256'h4189A45DE669556E506722ABD81E04DD3C52FBBB002B5D057123405147041041;
defparam prom_inst_2.INIT_RAM_3D = 256'h94C72F8A98172B734605A996692A4143DE2A8601546005188A9D420E7575CE86;
defparam prom_inst_2.INIT_RAM_3E = 256'h9582F501A7244AC82B1CD38D4A34A668AA80902ECE61A48253E1EB8CF0C032E5;
defparam prom_inst_2.INIT_RAM_3F = 256'hD3432441CC743BAA8BC8A2A284743C508F47D8D374B518C202739184733D8E95;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[29:0],prom_inst_3_dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 2;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hB00C60F2101C3F0F21CC721CCE0C70CFC413C413C41300D300D300D30FD34C3B;
defparam prom_inst_3.INIT_RAM_01 = 256'hC01D818F07D031960CB870C64509140BC2CB0002DC5CC0303044C5000600101C;
defparam prom_inst_3.INIT_RAM_02 = 256'h6D81E135C892711441B4F0CC1CC33C7B0CF020B2C05545455455455455155433;
defparam prom_inst_3.INIT_RAM_03 = 256'h2443F303C341C0C02D0361C300C3D804002D731C62C21C263F32FBECB32112C0;
defparam prom_inst_3.INIT_RAM_04 = 256'h5554000000000C1FFC0090FD0F00C3F00FD0FF00FC0FF0C3CC7830E01550004F;
defparam prom_inst_3.INIT_RAM_05 = 256'h360D0F0E1C30F3083090C70CB432F3CB0C0F61F3DC0FCB4343D081F31203CBC1;
defparam prom_inst_3.INIT_RAM_06 = 256'hF600073F18DB618BC3DFCCC040D0FD81F0F41F661F7F81FDCF4343C01320F184;
defparam prom_inst_3.INIT_RAM_07 = 256'hD0061C1044C02D00F3C074B1C0C0C0DFF0D614600D0030307FF2F0E618B387EC;
defparam prom_inst_3.INIT_RAM_08 = 256'h0871C7F610B3B01C32C0408CFFFF0BC7D80C0B1C30303030FD1C0FC0702C01C0;
defparam prom_inst_3.INIT_RAM_09 = 256'h4F343000D0300F3407F400CB1DCC1C1CFC61F7DF61C7600C71C21D4CD1C3C335;
defparam prom_inst_3.INIT_RAM_0A = 256'h00D01FD03431CCC7D040B0F20820830000E0E0CB32CF0F237D073433CCD304C3;
defparam prom_inst_3.INIT_RAM_0B = 256'h0303CC43031CC0C7430F3F57F3010C04D7F1D0F2C3EFF7BF0DEC04C000D0C3DD;
defparam prom_inst_3.INIT_RAM_0C = 256'h723FFFFD90C0343330C3C4394C0C70C303030D39F2731033FD3F00C725F30343;
defparam prom_inst_3.INIT_RAM_0D = 256'hCFB70C36398360B7C003FCC370DC370F33FD000183E063CBC62FFFC71CE4E81C;
defparam prom_inst_3.INIT_RAM_0E = 256'h4342CF35542594F646465A43C0B02CB1D08FD3FCFCBCBC022E4392CF03C82D3E;
defparam prom_inst_3.INIT_RAM_0F = 256'h1880C451451C93C0540C36596599143646464B0C8CCC2DAD12E41F1900951D94;
defparam prom_inst_3.INIT_RAM_10 = 256'h53C5305030850F13114053510C31D080BC30282CC0CC2CF0FDE320501E1E264E;
defparam prom_inst_3.INIT_RAM_11 = 256'h43CA581844451442C07F3D800DB7D856D6118461003C2C7F2CC2F55FC4451452;
defparam prom_inst_3.INIT_RAM_12 = 256'hC7F2C720054008CE0D0E40BC4034B3E4B2C7EC1F13CB6C361A41090614230BCC;
defparam prom_inst_3.INIT_RAM_13 = 256'h100310E1014010143C011630043111143D05433FFD0F438794073F2D84BDB503;
defparam prom_inst_3.INIT_RAM_14 = 256'hF1C7FC003800D90D01F107840F431E478767FE4E4E4E4E03D90D1F1079D0F433;
defparam prom_inst_3.INIT_RAM_15 = 256'h954B0F2C0041000F3FC78053D02D40FE4F2CF3FF170C0A36010F3C2D0C82CFD0;
defparam prom_inst_3.INIT_RAM_16 = 256'hCBFB4B82C202D101ED43C71D83DD0B502E03C70CB0C7FCC93CF02C4FA0363CBF;
defparam prom_inst_3.INIT_RAM_17 = 256'h171FCB92C7CBF3FCB888761091D87FC030330C00903F08503FD083C7A102F823;
defparam prom_inst_3.INIT_RAM_18 = 256'h47941B501E23FEB4740B6598B9C764BCFCBE47F3CBCFF30AC770E7F00C0CC000;
defparam prom_inst_3.INIT_RAM_19 = 256'hF8B401F3CDC0541009061D01C32CB30C33E5040743403FCF47C0054C0C023E10;
defparam prom_inst_3.INIT_RAM_1A = 256'h4F301503C0F7C06581047C00881043C0088104380B303010D82D40390C764024;
defparam prom_inst_3.INIT_RAM_1B = 256'hD051540C032E40F40C8000C1D03F0F0D2C34C03800430F1FC0443010CC0443CE;
defparam prom_inst_3.INIT_RAM_1C = 256'h32F372D4CECF1CBCC7D2CF933FC011014104BC10C92D42C10030100E0D050081;
defparam prom_inst_3.INIT_RAM_1D = 256'hFFF0FB02F2CFC3CBC8FF1FFC0C39DA00BF33FCCFF3C8CF81CF33CCF3073CC3C0;
defparam prom_inst_3.INIT_RAM_1E = 256'h7CF1CFC2F0C70C09003F4BFD01E470050CC407F37D9F3F3F2FFFCC7C3FFFF3F2;
defparam prom_inst_3.INIT_RAM_1F = 256'hD70140300332CB605C02F1FC0FCBC00C38B3E0E2F2C0CB0D38800D0FC72F073C;
defparam prom_inst_3.INIT_RAM_20 = 256'hB0C60F0CF3C342CF02FCC10207800C43CF041CD3340034003C3C307070D40240;
defparam prom_inst_3.INIT_RAM_21 = 256'hFCD00300FCF3CFCCF30F0DE9C10010CFC70390C7372C02C0D3CD0C0443C30000;
defparam prom_inst_3.INIT_RAM_22 = 256'hC07C7A1D9E71C3F878394BCB878B1C7A5C7F0C700C3320C02FC301C802CF0F33;
defparam prom_inst_3.INIT_RAM_23 = 256'hBF1FA830FC7CB06208FFF3C3F998CD60F9FC307000BB3FCB472702CB5C7A92D1;
defparam prom_inst_3.INIT_RAM_24 = 256'h27000BC3003B1F1C400CC907FBC7C3F30F1C710037240C7CCF2CF4040ED00FEC;
defparam prom_inst_3.INIT_RAM_25 = 256'h2C32F2CF03F02D0FC3C7C3F07F03FCB023C7873C43FCFFC00CD1C00377713C31;
defparam prom_inst_3.INIT_RAM_26 = 256'h00838F962F8300F4BC3C7D031964043CD1FF2C0CC0033C7CB0BC06464640CBFF;
defparam prom_inst_3.INIT_RAM_27 = 256'h0C11FCB02C82FC80013000A001402A00F002C013005C0F800581C509B8838080;
defparam prom_inst_3.INIT_RAM_28 = 256'h56107700B10B0FFC70CCC33B1C3B4078202C7F0FCB3D0D0C70FF1FC32DDF1E2E;
defparam prom_inst_3.INIT_RAM_29 = 256'h730040D81C3307F3FF2CFCF8791F30F3F1FFF3F0B12F1CBF00B80A05F694B614;
defparam prom_inst_3.INIT_RAM_2A = 256'h320BE1C31C1C3203F1CB2FCB3242C32070514236203D824CF333CD98C630F474;
defparam prom_inst_3.INIT_RAM_2B = 256'h5B6752614F644D320B3300B5802D02CF1CB1CBCBF1CB93A781A18E1024CB20BC;
defparam prom_inst_3.INIT_RAM_2C = 256'h7575D5757575575D75D575D72210030003215555555552221100333331028069;
defparam prom_inst_3.INIT_RAM_2D = 256'h5D575755D75D575775D55D57575755755755755755D5D5D5D755755D55775D5D;
defparam prom_inst_3.INIT_RAM_2E = 256'hD5755C5575D75D55D5777175D5755D575755755D5D5D57575D55D55D5D5D5D5D;
defparam prom_inst_3.INIT_RAM_2F = 256'h5D5D5D5C5C5C5D75D75D75D5D75D75D75D75D75D75D75EA75FAA575D5C55D715;
defparam prom_inst_3.INIT_RAM_30 = 256'h26666666665551323160000330203220230302023530022A1715715C5D75C5D7;
defparam prom_inst_3.INIT_RAM_31 = 256'hD4D4C5555555555541555555555408CCC084004C8448C40D5551301030031251;
defparam prom_inst_3.INIT_RAM_32 = 256'h800F10B1B3001CF031FF1F0F03C395C47B1001550554141551FD4100CF374704;
defparam prom_inst_3.INIT_RAM_33 = 256'h00F0D0305B30F583C081CE5C7370097371C6172DC21C718000001870F009C025;
defparam prom_inst_3.INIT_RAM_34 = 256'h31C303FDCCFF3C1C8720C70C0003F2F702718F07360B00F3DB2F0B247FCCBDCC;
defparam prom_inst_3.INIT_RAM_35 = 256'h15D80DB1DB3FC810363110F7731F3DCC3F3F0F73EDCBC76DCF3F3CD30D07C30C;
defparam prom_inst_3.INIT_RAM_36 = 256'h71871C572C0100701DC1170F60FF331457510C8558FF2C7F3C31F0C0C47C280E;
defparam prom_inst_3.INIT_RAM_37 = 256'h4C0C4C730347831D981E1CD1CDC18D621C300C373DC5872D86307018DB71C70B;
defparam prom_inst_3.INIT_RAM_38 = 256'h030032094F7601C0C0300C6000F000BFDFF73C9C1D0C2D4383F2DD038D5C1C1D;
defparam prom_inst_3.INIT_RAM_39 = 256'h03D583F2CB02FF0FD031CFF0F3CFEF63C3C70DCC0C3C3710B1F2DE79C0001851;
defparam prom_inst_3.INIT_RAM_3A = 256'hCF34F4403043CC3BF03F0C0B0C309063441E10B80D7770B8738DCF77F1CB2F0C;
defparam prom_inst_3.INIT_RAM_3B = 256'hFF423D8732C25C0C3033CB71C7009F63F1861CDBF2CC60B7E1FDC18F00C73031;
defparam prom_inst_3.INIT_RAM_3C = 256'h1C7CF013C014BC8FF001F7334B0C3F1F773CDF01010CE75F0F0FD5FC80C00000;
defparam prom_inst_3.INIT_RAM_3D = 256'h039C0918CB0B730F32C31430CF630C7CE363F1C0001DF1C7D8C7C01C1D9658FC;
defparam prom_inst_3.INIT_RAM_3E = 256'hD43091EF0BFCFCF1F3F03703D80D844D00C30CFC3FF73F0F1ACBC33B95400330;
defparam prom_inst_3.INIT_RAM_3F = 256'hD81EC30CB1C0C900027D87373C03E71C2D180B873331C744B0B50CB58E73DCCF;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[27:0],prom_inst_4_dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 4;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'hCCEE37DA3310221012042EAA5CB972EAD68B04ABCFB183BEFD7850A19236E28D;
defparam prom_inst_4.INIT_RAM_01 = 256'hEC7B0C224D603E1AD0C30C21E88305605E787F5D16DF3E2A778194D5BD8CAED8;
defparam prom_inst_4.INIT_RAM_02 = 256'h287337DE8BE38CE517ACECDAFEE78CF1062F6B0029C015EA24EB1DB00E0619A0;
defparam prom_inst_4.INIT_RAM_03 = 256'hDE8706A0C318AC73AD0E8AD0E48606A70DA984E60BA8809A70CA11A1DD85DFDD;
defparam prom_inst_4.INIT_RAM_04 = 256'hB9FFF6BBD38FC006400E4806A70EA1B30E0BA88B83ADCE19270CA13D9F10D3AD;
defparam prom_inst_4.INIT_RAM_05 = 256'hA0DF452F91ED0C2F18C70CA01371A053AD0E7CA03F06A380BA13AEAA70CA13D5;
defparam prom_inst_4.INIT_RAM_06 = 256'h06B5028DE3725D07AA6523D00E0923616DE88D906A87D181192AAE709A91270E;
defparam prom_inst_4.INIT_RAM_07 = 256'h6DDCF2830E2F60FA558C6F4A5B7E3DEA1B3D5918AD5BF86D02E51B128B07A18D;
defparam prom_inst_4.INIT_RAM_08 = 256'hBC6A6582E77790571CD5F4A5B7E3DEA11B3D3ADFE92A6E709A26270EA68CEE53;
defparam prom_inst_4.INIT_RAM_09 = 256'h426161FD5D62B70EA0000011B27B31F2CE587BE52ECA5231517F33532A1B189D;
defparam prom_inst_4.INIT_RAM_0A = 256'hD0F26D40012D3308E7B0A2B63E392A6E63E3207F5D0D452FE79012485F193187;
defparam prom_inst_4.INIT_RAM_0B = 256'hE0FAB2D09563E3363E333398ACD592D19BD17BD5391D2AA73E553E508299D296;
defparam prom_inst_4.INIT_RAM_0C = 256'h93D1E506B8F29D7DE2CEE0FA0829DA309022B9892D011A9D3363E513B21B72A4;
defparam prom_inst_4.INIT_RAM_0D = 256'h8A19FA3360FAF07E8D6082E3C27A98708297A7AA71EF03E384606E103A0324FD;
defparam prom_inst_4.INIT_RAM_0E = 256'hE5363E1D1383134275563E335A563EA6ADDD0FA711131A1E34AFEA536150A689;
defparam prom_inst_4.INIT_RAM_0F = 256'h11A352755814415504E81859151AFD5C8F632194DA1D3A308A546157B3616563;
defparam prom_inst_4.INIT_RAM_10 = 256'h219CDABD9511A163E99068F14C2A6A3EA42A4E8740A8E0FA888E800291785C15;
defparam prom_inst_4.INIT_RAM_11 = 256'h94D15885111A1D981121A84E0F219CD59F63E1906F5700A8B1ABD94D111D211F;
defparam prom_inst_4.INIT_RAM_12 = 256'h6A2E52AEEECAEED8DE502EDDECA92A8E7803AFD94D1AFDB578112113219FDAFD;
defparam prom_inst_4.INIT_RAM_13 = 256'hE91AADEAA5CB59F6DD8F7400E91C6D0AA57A02E9178D50AA7A03E14A6E54ABE8;
defparam prom_inst_4.INIT_RAM_14 = 256'h919BD503A3ADD699F35D5E27615AEEAFA4E1DA9E12A6E16A7E79A8E1DA5E7EA1;
defparam prom_inst_4.INIT_RAM_15 = 256'h11A1C5BE78CED35CD483BBCDB5311ABA4DCF35D681E975F706919747112B56DD;
defparam prom_inst_4.INIT_RAM_16 = 256'hDFF601FC903FD833EAD50CBF816A82B163E3E19ED55163E3E97D9963E968155E;
defparam prom_inst_4.INIT_RAM_17 = 256'hF5B92CF5B606E57A111AFD5973697736508E0FA36311127FCFFDAFD3ADA6289D;
defparam prom_inst_4.INIT_RAM_18 = 256'h3E8681E484E485E26562180EDDD87F98EDD587FF97AEDD60E2F65631CF87B92C;
defparam prom_inst_4.INIT_RAM_19 = 256'h3709AB03CFA981F0BAB09A550C2F69A86E64270CA70F2A9B169111506FF61688;
defparam prom_inst_4.INIT_RAM_1A = 256'h6B0B2900D2195D51950DA333506F5531581F53168F4115531CF8906533E6CA8A;
defparam prom_inst_4.INIT_RAM_1B = 256'h8CEE7CB53B11E5D55730EA591112981607112F711429311F7913B2331331A0F0;
defparam prom_inst_4.INIT_RAM_1C = 256'h30E75A619222E70EA00363E33E8E4039E803E780FAFB0DAB9E0BA50E210329FE;
defparam prom_inst_4.INIT_RAM_1D = 256'hF06B0D29CD789BB25D0D1BAD5303131200B1970EA310823393DF3031106F3792;
defparam prom_inst_4.INIT_RAM_1E = 256'h227968948469D40FAB0D4D19BAD7D2F53363E163EF70813233BBB99BE08A73A0;
defparam prom_inst_4.INIT_RAM_1F = 256'h9DAA37FF06AC637ACF3D06AB00A86D9ADD079001B0DA97174D0F25F903AB9197;
defparam prom_inst_4.INIT_RAM_20 = 256'h19AD85DFDD9236E015C302A59156D906F81176590EAB19AC3E50FA580155CD71;
defparam prom_inst_4.INIT_RAM_21 = 256'hB33D8C2E40838A687CE3FE5026B912333750318FD919EDF58AD63E18FD53E5AB;
defparam prom_inst_4.INIT_RAM_22 = 256'h728313CDE3ADA85494D9AD85D3923EE0E1032F06193D0F23E11203A5E0318AD9;
defparam prom_inst_4.INIT_RAM_23 = 256'h871FB03AB051500A500106201A58115F92AAE191B306278F39F6FF06AB00A51E;
defparam prom_inst_4.INIT_RAM_24 = 256'hB39906E1082B03E9592D3E9BAFB0DAB168906FF9BD403E333E38FB0BAB09A9A2;
defparam prom_inst_4.INIT_RAM_25 = 256'hAD4B90906EB5EB6B84D11955511109053F31890F06AD48363E36F59F1A8FB08A;
defparam prom_inst_4.INIT_RAM_26 = 256'h9196D96DB04A59DD39ED187D92ACE6511A5EA4D34FD311A55893B09031198D06;
defparam prom_inst_4.INIT_RAM_27 = 256'h20FBEB6B03A910629750F06AEB9050B95DB11AA4D88332A8DCF63E3E31843533;
defparam prom_inst_4.INIT_RAM_28 = 256'h7539F37DCF5BCD8F78431304ABFD87D1E9A63E3EAAA7D578197E7F97D5781903;
defparam prom_inst_4.INIT_RAM_29 = 256'h06863635118FD50E18288E55EF3FAFDA8B0D3704A48DC1F87DB551A3D38BFD58;
defparam prom_inst_4.INIT_RAM_2A = 256'h1EF006ED5A91319FBCDCF589EFE5EAA54A2DEBB80A51AFD8439ED19EDF8ADD49;
defparam prom_inst_4.INIT_RAM_2B = 256'h63BED78303D042BFD193972AE935119FB9011E5DE532695F63E3F78AA7D9387B;
defparam prom_inst_4.INIT_RAM_2C = 256'h8363E11022FF15B0D10C21E9B7BEA2B5D37D718CF072042BCD97A1BAFD537D70;
defparam prom_inst_4.INIT_RAM_2D = 256'hA57833AD87EE80EDB5D07ABED3AD10EFFD0C2B553A8A1FB35363E5DBD1FDA9A1;
defparam prom_inst_4.INIT_RAM_2E = 256'h73E88A532F670DBC237E601F5F6B4C5E4444BBBB80BE0D3827E385306A31D407;
defparam prom_inst_4.INIT_RAM_2F = 256'hEA3D537D24D90929090F332A09AB3A81187D991EA2F53D450BCD551B0D681B72;
defparam prom_inst_4.INIT_RAM_30 = 256'h001BDC112771FAA3D37D787E53F1F28269118D80F24D3A09AB04A24DA21D24D3;
defparam prom_inst_4.INIT_RAM_31 = 256'h99118D092A02CDD037E9CD31026F25D3604A70B38DC25D70703625D36B11A23D;
defparam prom_inst_4.INIT_RAM_32 = 256'h38D921BCDCF5B2D783EAFD0D4122826D8080725D36CE2A8387D1DDA83504A87D;
defparam prom_inst_4.INIT_RAM_33 = 256'hE9D5E3120C300EE7A5E3E2E58C8963E3EAA0655A0E2F5B1C870EA8811ABBFA4D;
defparam prom_inst_4.INIT_RAM_34 = 256'h0E4EE3832E880AE484E00ED85E08EE3EB788EBEDEA5783EE4A1E3E7E9D7FF3AD;
defparam prom_inst_4.INIT_RAM_35 = 256'h45D715683E3E585C31E00EE3EE68706AA0CE083E88EE3E7850EC72C306FEC570;
defparam prom_inst_4.INIT_RAM_36 = 256'h1137D550811572468E70EE68D6E0878D5086CBA1BA34711846830E30E30E0BED;
defparam prom_inst_4.INIT_RAM_37 = 256'h9D68D32789F06963E30E5551B17972CE58BE0E2D877B187DFED06AEA29E18355;
defparam prom_inst_4.INIT_RAM_38 = 256'h40E76111A8ADA8D50E111A551A4D37D59811E9D51E1E19319DD30ECCB2113ADE;
defparam prom_inst_4.INIT_RAM_39 = 256'hFD51BED5363E3390E92BCDB0C2B10EFD488BC540AA0A2913A4BE7A5783ADD3A5;
defparam prom_inst_4.INIT_RAM_3A = 256'hF2A8E4EB2453E915B8737277AFA0AEE80634D0671A037ECFE53ADEE07A3AD0EF;
defparam prom_inst_4.INIT_RAM_3B = 256'hEF5A8EC8BEF8A8EF3A5EF5A3EFAA4EFDA9EF83EF0ACEF6A1E06281E180EF0ADE;
defparam prom_inst_4.INIT_RAM_3C = 256'h91805B0BE4328F1C513ADFEA7EFFC51F34D573FF15950533AD487EE530ED1101;
defparam prom_inst_4.INIT_RAM_3D = 256'h34DFADF68069105433AD734D87E93AD1E305F1D3AD987E3AD1E87EEC310EDB5D;
defparam prom_inst_4.INIT_RAM_3E = 256'h6FB54C048138FE953837BE380A77ED55FD15B3ADF8458EE08BEF0ADEA88EFDA7;
defparam prom_inst_4.INIT_RAM_3F = 256'h2433EA9311A835378B07AC3A110EDB5D93053AD8EB5878FD333AD71198D3D490;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[27:0],prom_inst_5_dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 4;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'hC2F723C13CC4E2E4E34E214CB7E19C15C02E4E2E2CE12EE14C12D0011AC21032;
defparam prom_inst_5.INIT_RAM_01 = 256'hFCD249308C022F4CC27C49303E1F21F29FDCB10C0115C1CDD02E09CE217CCF17;
defparam prom_inst_5.INIT_RAM_02 = 256'h32EE23C523F522FE23CBF2BCBF7C12CE4A33E74221302E14D0F20C126F2F26C2;
defparam prom_inst_5.INIT_RAM_03 = 256'h03CB4A327CE2ACB02C232AC2FDB84A34493018F8493022EFB4934224CC26C0BC;
defparam prom_inst_5.INIT_RAM_04 = 256'h22C57E21C212F31D332FDB4A3449322C7F493024102C2321FB4934DCCA4DC02C;
defparam prom_inst_5.INIT_RAM_05 = 256'h30044453C4BC493A0FFB49328CDEF2002C234303824A30149325C14FB4934DCE;
defparam prom_inst_5.INIT_RAM_06 = 256'h032F1020F2703C4A2F0E09C2274A32D4DC722CC4E22AC272C1AC21B4A319CB4D;
defparam prom_inst_5.INIT_RAM_07 = 256'h20C2C01E4D3AF4F2E012310CC2B721BDC1BCECE2ACE3C26CC2FC2D02124A20FC;
defparam prom_inst_5.INIT_RAM_08 = 256'h22031022F45D12FE4DCD10CC2B721BDCD1BC02C331AC01B4A329CB4D3222F7DE;
defparam prom_inst_5.INIT_RAM_09 = 256'hC282B4DCD19CEB4D300000D2FCD2E27C2F02D206D06DC240FFD13CDE252EF26C;
defparam prom_inst_5.INIT_RAM_0A = 256'hC4D220C00122CE28FDE4D2E52521AC01B27212B10C006676666267774326CE2A;
defparam prom_inst_5.INIT_RAM_0B = 256'hF4A30DC66E525E242422222100CE0CCE0CCE00CEE0BC2EFB27DF27D4E2F19C13;
defparam prom_inst_5.INIT_RAM_0C = 256'h16C00D0122C2BCD11C2F74D24E2F11C664A2E020CC9CE03CE2525DE727EE0BC0;
defparam prom_inst_5.INIT_RAM_0D = 256'h19228CB0D4A35D0FDCD4D272ECB7E1D4D219D5BA10F030F13DD017C4F24F229C;
defparam prom_inst_5.INIT_RAM_0E = 256'h4C2424412032F2CEBFC42422CFC4240FC3334A3B4222ED5F2DC7F7C240CDB571;
defparam prom_inst_5.INIT_RAM_0F = 256'h42229CEE2B2601DCD6F7E12E0ED07CDE1711F00AC0BC23C4D2C200C440CF0C42;
defparam prom_inst_5.INIT_RAM_10 = 256'h2E0FC0DCCC422D42400001B227D0FC0F727C0F7526C0F4A3220F74B37CC1280E;
defparam prom_inst_5.INIT_RAM_11 = 256'h0ACED11B2DC0BCD1422ED20F4A3F0FCCE6627C0004C04B31A20DC0BCDC412E41;
defparam prom_inst_5.INIT_RAM_12 = 256'h6C2F23CCF06C2FE2CF24D13C06D1AC21D0AC0CC0ACE0CCEEE1422E422E0BC0CC;
defparam prom_inst_5.INIT_RAM_13 = 256'hFCE09C14CB7EE2C20C2CD12CFCE06C4E2ED02CFCE2FCE493D02CF49C2F2CCCF2;
defparam prom_inst_5.INIT_RAM_14 = 256'hCE07CE4F223C71C2C23C24DDD45CBF22CCF09CCF03CCF47CCF2CCCF49CCF2FCC;
defparam prom_inst_5.INIT_RAM_15 = 256'h1E0BDE1F030F7E22C11EE21CEEE422E0FC2C23C134F7DC4000CE0FCE422EE20C;
defparam prom_inst_5.INIT_RAM_16 = 256'hC9FCAC8306C3E202B011D3BAD0D7CB7E42425D2DCFCD424272DCE66240100D23;
defparam prom_inst_5.INIT_RAM_17 = 256'h6A7CB76B7024FC2F0DF07CCCB0DC3B0D030F4A324CC42262762707C23C511108;
defparam prom_inst_5.INIT_RAM_18 = 256'h2F01C2F1C2F1C2F01D251F313CF3D40313C03D4A19D13C44A3AFC2002CCD2CA7;
defparam prom_inst_5.INIT_RAM_19 = 256'h102B1021B6112ED4F2E4F2DE4D3A2EC2D726CB4D3D4A37C2E51402E0157E4D7C;
defparam prom_inst_5.INIT_RAM_1A = 256'h324F2664F2E15CEC0E4F2000C004CEEF32DD24132D2F1DFEE7D1102E1132CCB1;
defparam prom_inst_5.INIT_RAM_1B = 256'h22F753EEEEFC14CCD5E4A2ECE42212202E42266C423CEFF55CE1E727D27DF2D0;
defparam prom_inst_5.INIT_RAM_1C = 256'hC1129C9F1AC11B4A3E22525223B7022B7022B224A3DE4F2E134F2D4A2E4F22CE;
defparam prom_inst_5.INIT_RAM_1D = 256'hD0324F216CC31E44FE23F0ACF27270C03000714A3274D22216C42727F015271A;
defparam prom_inst_5.INIT_RAM_1E = 256'hCEB2022030D2444A3E2443F10AC23DDFE2525E1274433F272722E02E54D250F2;
defparam prom_inst_5.INIT_RAM_1F = 256'hAC09C6A64A306C6976974D2E4A22EC2DC02E3002E4F2CDE2DC4A3EAC4F2E0C02;
defparam prom_inst_5.INIT_RAM_20 = 256'h02DC26C0BC1AC11CEB724A2ECE28C00041A20EEE482EF2DC0FF4A3E092E22CD4;
defparam prom_inst_5.INIT_RAM_21 = 256'hE2E17C2FF2B02B02B072F0E5202CE72727E4D22BCCD2CC6E25C424E2BCE27C22;
defparam prom_inst_5.INIT_RAM_22 = 256'hBF1020C0F02C0C110CC2DC26C21AC11C7E4B2D4D10DC4A3034224B2D34D125C7;
defparam prom_inst_5.INIT_RAM_23 = 256'h2F0DE4B2E4B2E4A2E0024D24B2C2C0FB1AC11FCFE24D203D20F0424D2E4A2FF0;
defparam prom_inst_5.INIT_RAM_24 = 256'hE200004E4D2E20F0E0CC2726CDE4F2ECE11015A24C020F222712DE4F2E4F224C;
defparam prom_inst_5.INIT_RAM_25 = 256'h24425500262E4242CB7EDCCDEFFCD66EEDEED66D4D244C25252BAC230D2DE4D2;
defparam prom_inst_5.INIT_RAM_26 = 256'h422CC2CCE4D2E2DCE2DCD25C1AD118E422E70FCE29CE422EC2EC266727E15C4D;
defparam prom_inst_5.INIT_RAM_27 = 256'h2CD242424B2CE4D20402D4D24155DCE2FCE4220FCF11010C22642427EE28CEE2;
defparam prom_inst_5.INIT_RAM_28 = 256'hEEE2C23C2CD21C2CD28CC74D221C25C03C1525214C20CC2F0CB75A2DCC2F0C4B;
defparam prom_inst_5.INIT_RAM_29 = 256'h0066242EEC2BCC001703B7EE34EA2DCC1F21274D2D211F525C7FFD21C0121C02;
defparam prom_inst_5.INIT_RAM_2A = 256'h974D00B3C260EF2C21C2C022FF1C14C002EC7EC191DD2DC28C2DCD2CC625C440;
defparam prom_inst_5.INIT_RAM_2B = 256'h9C20C2FC49C49321C4DC19C7FC4CDC2CEC7EC06C7CE741E6627252FC20CC4D4B;
defparam prom_inst_5.INIT_RAM_2C = 256'h72424DE4A2FF2C11CC49303C7D214C20C23CD012C49349321CCB7EE07CE23CD4;
defparam prom_inst_5.INIT_RAM_2D = 256'h2EF1202CCB7B12FC27C4A227C02CE230AC4E2ECEE11DCDEEC2424C19C4DC11CB;
defparam prom_inst_5.INIT_RAM_2E = 256'hB272DC1007EF212AF2B71525E7D02C9F1111000002FF32CC0B72C10009CE444A;
defparam prom_inst_5.INIT_RAM_2F = 256'h321CE23C08CC4F266F2D10014F2EE1E2C2AC12214DDEE550312CCCD11CC1E2BF;
defparam prom_inst_5.INIT_RAM_30 = 256'h00214C4226BF6121C23C02B7F220A02BDCE0FCF2D06C114F2E4A206C106C06CD;
defparam prom_inst_5.INIT_RAM_31 = 256'h1220FC4F2E102CE22B716C722A9503C004A232B021103CF1F2DD03C00E42209C;
defparam prom_inst_5.INIT_RAM_32 = 256'h23CC1D21C2CD20C2FC707C00444A109CF1F2B03C0033311C2AC3BC1ECE4A22AC;
defparam prom_inst_5.INIT_RAM_33 = 256'h24C234EF10022F21C2F2700E5116624214CB4DFB4D3AEED02B4D301422E3C0FC;
defparam prom_inst_5.INIT_RAM_34 = 256'h232F70320F7C22F122FD2BB22F422F272E2032F2FC0322F21C2F27524C55A02C;
defparam prom_inst_5.INIT_RAM_35 = 256'h5D291DF22F27220020092232F7E154F7122FF22F122F2742000158121CAF1002;
defparam prom_inst_5.INIT_RAM_36 = 256'hCD23CDC52FE0580C0302FF022D712B71120E127DEC214DDD0D72CB2CB2CBC5F5;
defparam prom_inst_5.INIT_RAM_37 = 256'h4C0120CB715016624297DFEEECD19C2F023F4D3023D2E2AC0BC8F714D1F874EC;
defparam prom_inst_5.INIT_RAM_38 = 256'h02349F4222AC26CC004422ECC0FC23CCE2FE24C0F30026CE2DCE2FD2CCFE02C2;
defparam prom_inst_5.INIT_RAM_39 = 256'hACEE27CC242422661DD12CE4E2EEC14C01CE3AB4E2493CF02C23B7FF102C2DC0;
defparam prom_inst_5.INIT_RAM_3A = 256'h2DCDF12BC11E292EE158080075030F033D08C014EF22B70F0E02C034A202C230;
defparam prom_inst_5.INIT_RAM_3B = 256'hF27C1F121F27C2F2EC1F26C1F24C1F27C1F322F24C1F2FC2F2D033F42FF2ECDF;
defparam prom_inst_5.INIT_RAM_3C = 256'hCFE21E2B702032ADFF02C23CB725DFF508CF3E252ECF21202C0CB726C2FCDCC1;
defparam prom_inst_5.INIT_RAM_3D = 256'h08C20CF1403CF210202C708CCB7C02C23F212AC02C02B702C23CB727CC2FC27C;
defparam prom_inst_5.INIT_RAM_3E = 256'h26EC009C1F03FF7FF12727209C3B70ED2710202C12000312C1F2EC0F020F27CB;
defparam prom_inst_5.INIT_RAM_3F = 256'hB4CCD11CDC19CF23C24A23A7DC2FC27CCF2102C0320CB727C202C7FC15C24410;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[23:0],prom_inst_6_dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_2),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 8;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'h5AC335FBC335C2C33455C334ABC331D1C331C0C332DAC33274C3329BC3325EC3;
defparam prom_inst_6.INIT_RAM_01 = 256'h351CC36FCBE4DB35A0C335BBC33799C3377BC331F7C33739C3338EC33680C336;
defparam prom_inst_6.INIT_RAM_02 = 256'h7A797877767574737271706F6E6D6C6B6A6968676665646362614037B5C3D318;
defparam prom_inst_6.INIT_RAM_03 = 256'h05DC212009080A5B011F0D2F2E2D2C3B3A39383736353433323130C9B737EA3A;
defparam prom_inst_6.INIT_RAM_04 = 256'h5A595857565554535251504F4E4D4C4B4A49484746454443424160C9AF41FF22;
defparam prom_inst_6.INIT_RAM_05 = 256'h21013E2019181A1B011F0D3F3E3D3C2B2A29282726252423222100AAAAC9AF77;
defparam prom_inst_6.INIT_RAM_06 = 256'h5A595857565554535251504F4E4D4C4B4A49484746454443424140DB18AE4019;
defparam prom_inst_6.INIT_RAM_07 = 256'hA6E1282009080A5B011F0D2F2E2D2C3B3A39383736353433323130C9AF01D9CD;
defparam prom_inst_6.INIT_RAM_08 = 256'h5A595857565554535251504F4E4D4C4B4A49484746454443424160C9EFC001FE;
defparam prom_inst_6.INIT_RAM_09 = 256'h41FD3A2019181A1B011F0D3F3E3D3C2B2A29282726252423222100C901CB2314;
defparam prom_inst_6.INIT_RAM_0A = 256'h3A393837363534333231302F2E2D2C2B2A29282726252423222120C941FE3A6F;
defparam prom_inst_6.INIT_RAM_0B = 256'h5A595857565554535251504F4E4D4C4B4A494847464544434241403F3E3D3C3B;
defparam prom_inst_6.INIT_RAM_0C = 256'h7A797877767574737271706F6E6D6C6B6A696867666564636261405F5E5D5C5B;
defparam prom_inst_6.INIT_RAM_0D = 256'h2CA521C9FE10780631F3CDFE100D06FFD3023EFE100D06FFD3013E7F7E7D7C7B;
defparam prom_inst_6.INIT_RAM_0E = 256'hCD3C3E53ED202011ECDBEBE5C5E3EBC9FB31EDCDFDE642103AFFDBE0D342133A;
defparam prom_inst_6.INIT_RAM_0F = 256'h2B01CD0253C223D67EC9FFD3AFC9ECD342103202F642103A0060C37D000131E8;
defparam prom_inst_6.INIT_RAM_10 = 256'h78187A3C3F320AEE3C3F3A08204212325FE63C42123AFB103220CD0806C92CCF;
defparam prom_inst_6.INIT_RAM_11 = 256'h1812CB17C1FFDBFE10980631F3CDFE106E06335CC3F628028DCD083817FFDBC5;
defparam prom_inst_6.INIT_RAM_12 = 256'h21E5F318FE109A06C9F1C1D1F3200D31A5CD0A3002CB31A5CD57080ED5C5F5B2;
defparam prom_inst_6.INIT_RAM_13 = 256'hCD00164006420E22320321E523183241CDA53EFB103241CDAF5306420C223241;
defparam prom_inst_6.INIT_RAM_14 = 256'h2232BA21E5C9D1C1E17C3C3E222A2A21F820A5FE7A3220CDF710F520B77A3220;
defparam prom_inst_6.INIT_RAM_15 = 256'h3ECD4FD5C5F507184FD5C5F5E318A53E32B4CD7F3EF91032B4CD553E0006420C;
defparam prom_inst_6.INIT_RAM_16 = 256'h0E2232CA21E5320AC3F810337CCD3350CD08063350CD8A18FB103335CD080633;
defparam prom_inst_6.INIT_RAM_17 = 256'h3350CD3350CD4006000021F210F2303EFEF6380FFE793350CD8006E0D3013E42;
defparam prom_inst_6.INIT_RAM_18 = 256'h023ED720BD0A28BC403EE4102C0318E9102405380DFE44ED0230917A3350CD51;
defparam prom_inst_6.INIT_RAM_19 = 256'h2F110318121711053001CB3290C3F5207FFE7A337CCD3350CD00163350CDE0D3;
defparam prom_inst_6.INIT_RAM_1A = 256'h224B4221F3F82804E638403A0C000EFBC9FFD3013EFD201DFFD3023EFD20152B;
defparam prom_inst_6.INIT_RAM_1B = 256'hCB22FE79C9FBF1C9F1F10320BB01E6FFDB4F81063E001E0218011E4203C33C3E;
defparam prom_inst_6.INIT_RAM_1C = 256'hC300C401500021C0FEFEC4DBC5D3033E1318C93C3E32443ED83EFE03380FFE12;
defparam prom_inst_6.INIT_RAM_1D = 256'h0A00164036213801014224321F3E022846CB25CB082866CB384021FF3E003417;
defparam prom_inst_6.INIT_RAM_1E = 256'h222342012AE5307DC342012262ED0820A6313DCD33BFF23120CD3220A373AE5F;
defparam prom_inst_6.INIT_RAM_1F = 256'h0060CD05C401C55FAB1841FF22962E42012212AF30A1DAD152ED41FF5BED4201;
defparam prom_inst_6.INIT_RAM_20 = 256'h803A00005000C3B2EDFA18140A380F7B571717177A41FD327D41FE32C8A30AC1;
defparam prom_inst_6.INIT_RAM_21 = 256'hBDCAB74730A1CA1AFE7E1900165A304521FACB0228B740193AF2CB022803E638;
defparam prom_inst_6.INIT_RAM_22 = 256'hECD320F6E4D3407D3156ED3390C337AFC230FDC378BE1F3E04202AFE42242130;
defparam prom_inst_6.INIT_RAM_23 = 256'hF921B0ED004C0140001136AA21F0D30B3EE0D3043E3518CDF0D3D03EF4D3813E;
defparam prom_inst_6.INIT_RAM_24 = 256'hF4D3813E0B00000137AFCA3CF0DB344FCD028DCD01C9CDB0ED00400141E51136;
defparam prom_inst_6.INIT_RAM_25 = 256'h21F120B178F4D3813E0B11204FCBF0DB000001051EF02857CBF0DB37AFCAB178;
defparam prom_inst_6.INIT_RAM_26 = 256'h00F301E4D3803E404932C33E404A22350221F4D3813EE3201DE418021BCD0277;
defparam prom_inst_6.INIT_RAM_27 = 256'hC3A2EDF4D340F6813EA2ED34EECA02E6F0DB3518CDF0D3803EF2D3013E430021;
defparam prom_inst_6.INIT_RAM_28 = 256'hDB4049C2C900C1C5B2184300CA1CE6E1F0DB3518CD40492245ED21E4D3AF34F7;
defparam prom_inst_6.INIT_RAM_29 = 256'h2035401A211C20B7401C3A2228B740223AECDBD5359111FF0000C3FA286FCBE4;
defparam prom_inst_6.INIT_RAM_2A = 256'h11231E36C03542162177203E021840233A052840202A7701EE01E67E23073616;
defparam prom_inst_6.INIT_RAM_2B = 256'h237E2B06301EFE7ED0BE1A5F833D2B7E233423F710132377C0961A3403060266;
defparam prom_inst_6.INIT_RAM_2C = 256'h3C3521C01EFE42163AC847CB42103AC9342B2B0136D80DD67E34230136C803E6;
defparam prom_inst_6.INIT_RAM_2D = 256'h2F0E421C11EC182371C8052377233AC6FB300AD6342F361B1A03063A0E421911;
defparam prom_inst_6.INIT_RAM_2E = 256'h403DD21F4046D21FE535F121E5FDE5DDE5D5C53369D21F3365D21FE0DBF5E318;
defparam prom_inst_6.INIT_RAM_2F = 256'hFFFEEADBF3C9FBF1C1D1E1E1DDE1FDE14043D21F4040D21F4209D21F4206D21F;
defparam prom_inst_6.INIT_RAM_30 = 256'hFD0428B7057EDD3644CD41E521FDEAD32A28B7047EDDE9D3037EDDE8D3AF3828;
defparam prom_inst_6.INIT_RAM_31 = 256'hEDE80E0406AFC9FBE8DBD604CBFDCE04CBFD0428B741ED21FDD604CBFDCE04CB;
defparam prom_inst_6.INIT_RAM_32 = 256'hDDAF41E521DDDC18FB10230036030641F021FB10230036030641E821FB100C79;
defparam prom_inst_6.INIT_RAM_33 = 256'hC90377DDEBDB4203C3F028028DCDC84E04CBDD0D207FCBEADBC85604CBDD0377;
defparam prom_inst_6.INIT_RAM_34 = 256'hB7037EDD4203C3F028028DCDC84E04CBDD0D2077CBEADBC85604CBDD41ED21DD;
defparam prom_inst_6.INIT_RAM_35 = 256'h013018C30000C90000C925D9C31C90C31D78C31C96C3C9000336DDEBD3790120;
defparam prom_inst_6.INIT_RAM_36 = 256'h00C9AF0000C75000C352FF00014303C20600B0003C0004730700000701003024;
defparam prom_inst_6.INIT_RAM_37 = 256'h52000000301E010000000000C73529C335FAC335FAC335FAC3AAAAAAAAAAAAAA;
defparam prom_inst_6.INIT_RAM_38 = 256'h35FAC335FAC3022EC30000FFFF00004E52FF6C55301B024F5200000030210249;
defparam prom_inst_6.INIT_RAM_39 = 256'h032052FE037EDDFF000000003739020000000000001E0000043C033832033241;
defparam prom_inst_6.INIT_RAM_3A = 256'h6C21C9B0ED000301C0E1EB375ECD067EDD032052FE057EDDE5C0375ECD047EDD;
defparam prom_inst_6.INIT_RAM_3B = 256'h3A0A2022FE41ED4F41E549402550401D4440154BC96F66237EC0B1ED000F0137;
defparam prom_inst_6.INIT_RAM_3C = 256'h2857CD113EE5D706A3C31706A8DA1F409F3A06AAC23AFE223E409F3201EE409F;
defparam prom_inst_6.INIT_RAM_3D = 256'hCD021BCD37F62137D7CDFB0075C337B5CD2884C335A0CD23203635BBCD40D42A;
defparam prom_inst_6.INIT_RAM_3E = 256'h223030210033C30D3E421132AFE2204CFE052848FEF10033CDF50E280DFE0049;
defparam prom_inst_6.INIT_RAM_3F = 256'hAAAA03203F737361430EE618021BCD020221021BCD01FFFFAAAAAA022EC34177;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[13]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[12]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(prom_inst_4_dout[0]),
  .I1(prom_inst_6_dout[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_5 (
  .O(dout[0]),
  .I0(prom_inst_0_dout[0]),
  .I1(mux_o_4),
  .S0(dff_q_0)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(prom_inst_4_dout[1]),
  .I1(prom_inst_6_dout[1]),
  .S0(dff_q_1)
);
MUX2 mux_inst_11 (
  .O(dout[1]),
  .I0(prom_inst_0_dout[1]),
  .I1(mux_o_10),
  .S0(dff_q_0)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(prom_inst_4_dout[2]),
  .I1(prom_inst_6_dout[2]),
  .S0(dff_q_1)
);
MUX2 mux_inst_17 (
  .O(dout[2]),
  .I0(prom_inst_1_dout[2]),
  .I1(mux_o_16),
  .S0(dff_q_0)
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(prom_inst_4_dout[3]),
  .I1(prom_inst_6_dout[3]),
  .S0(dff_q_1)
);
MUX2 mux_inst_23 (
  .O(dout[3]),
  .I0(prom_inst_1_dout[3]),
  .I1(mux_o_22),
  .S0(dff_q_0)
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(prom_inst_5_dout[4]),
  .I1(prom_inst_6_dout[4]),
  .S0(dff_q_1)
);
MUX2 mux_inst_29 (
  .O(dout[4]),
  .I0(prom_inst_2_dout[4]),
  .I1(mux_o_28),
  .S0(dff_q_0)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(prom_inst_5_dout[5]),
  .I1(prom_inst_6_dout[5]),
  .S0(dff_q_1)
);
MUX2 mux_inst_35 (
  .O(dout[5]),
  .I0(prom_inst_2_dout[5]),
  .I1(mux_o_34),
  .S0(dff_q_0)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(prom_inst_5_dout[6]),
  .I1(prom_inst_6_dout[6]),
  .S0(dff_q_1)
);
MUX2 mux_inst_41 (
  .O(dout[6]),
  .I0(prom_inst_3_dout[6]),
  .I1(mux_o_40),
  .S0(dff_q_0)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(prom_inst_5_dout[7]),
  .I1(prom_inst_6_dout[7]),
  .S0(dff_q_1)
);
MUX2 mux_inst_47 (
  .O(dout[7]),
  .I0(prom_inst_3_dout[7]),
  .I1(mux_o_46),
  .S0(dff_q_0)
);
endmodule //Gowin_pROM_M3
