//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-4 Education
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Fri Jun 07 22:50:11 2024

module blk_mem_gen_0 (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [7:0] douta;
output [7:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [11:0] ada;
input [7:0] dina;
input [11:0] adb;
input [7:0] dinb;

wire [11:0] dpb_inst_0_douta_w;
wire [11:0] dpb_inst_0_doutb_w;
wire [11:0] dpb_inst_1_douta_w;
wire [11:0] dpb_inst_1_doutb_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[11:0],douta[3:0]}),
    .DOB({dpb_inst_0_doutb_w[11:0],doutb[3:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[3:0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b0;
defparam dpb_inst_0.READ_MODE1 = 1'b0;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 4;
defparam dpb_inst_0.BIT_WIDTH_1 = 4;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'h3F009023008E30F300B830C300B4309300253063002930330085300307869463;
defparam dpb_inst_0.INIT_RAM_01 = 256'h069460303C3F005C54FDA83053999E88E00110F56D90D332E3E0010B176C30E4;
defparam dpb_inst_0.INIT_RAM_02 = 256'h00000000000000000390EF932560DF204FF29C3C0BAC3F00038D43FD81096181;
defparam dpb_inst_0.INIT_RAM_03 = 256'h0513D4060510D03109105126D430E26D430EC227B80A80B931DE0F1F6030E6D0;
defparam dpb_inst_0.INIT_RAM_04 = 256'h001D00EC88EC84871AD807E7810D506E09A681F1E26586E07278F461E57FF10D;
defparam dpb_inst_0.INIT_RAM_05 = 256'h281BD50706A1A47F7DC5C86B6375E073FFFF63E9F06231748CAA3E68700170C1;
defparam dpb_inst_0.INIT_RAM_06 = 256'h003C30E43F985680AF431B8705A0420821E401126D55A2DF411001431E780FBD;
defparam dpb_inst_0.INIT_RAM_07 = 256'h911F0ED903330E3EA600190EE825CD062B0F301001052C11C0707A682E0F162E;
defparam dpb_inst_0.INIT_RAM_08 = 256'h39F0D0E135D4001431E001BD803A8EDEE6301D0704A90D3D473F1C010E90512D;
defparam dpb_inst_0.INIT_RAM_09 = 256'hF3935332B272DA87781540C8CDA0C73AF3AD4363E488833287E7C6A95E07E535;
defparam dpb_inst_0.INIT_RAM_0A = 256'hE5149434BFF7D7177707D4910FE4969515A4500FE49494045474D47373531373;
defparam dpb_inst_0.INIT_RAM_0B = 256'h65C767D4910FE6B5C636D5A634500FE5F5C45FF7D78704B4310FE6056434B00F;
defparam dpb_inst_0.INIT_RAM_0C = 256'hD10FE6D5A5F00FE5049425D5047FF7771717D10FE6D566300FE5049425847FF7;
defparam dpb_inst_0.INIT_RAM_0D = 256'hF00FE5149425D5047FF7D787071717D10FE60566300FE5149425847FF7778717;
defparam dpb_inst_0.INIT_RAM_0E = 256'h0FE5D50575D575DFF7210FE655F00FE5E42504757FF7D787078717D10FE60565;
defparam dpb_inst_0.INIT_RAM_0F = 256'hD505C4547FF7B7A737B10FE61686A00FE5D50575D52FF7B7A757B10FE61685D0;
defparam dpb_inst_0.INIT_RAM_10 = 256'h752FF5752FF7778717D5C767D4910FE6D5610FE5F5C636D5A634500FE5049425;
defparam dpb_inst_0.INIT_RAM_11 = 256'h17B5C727A7110FE6E596710FE5D665C694500FE53565700FE595450454700FF5;
defparam dpb_inst_0.INIT_RAM_12 = 256'h41FC00584FF8A5C7D718B10FE635C6D6D4500FE5B5C454CFF8C59885D10FE777;
defparam dpb_inst_0.INIT_RAM_13 = 256'h04FE039004FF20045E3210000569240EF04E5F6004FE031700571D90DF2007E9;
defparam dpb_inst_0.INIT_RAM_14 = 256'h3940421800900FC6034E548509E1D0FF400D04541FC052047E13005C21C91610;
defparam dpb_inst_0.INIT_RAM_15 = 256'h323001414043FC00E9171092404E102FF40053FC30094152052105F90E58700B;
defparam dpb_inst_0.INIT_RAM_16 = 256'h315C0004E103B39408349730E5520318002584FE1053502F00C02F2250B55300;
defparam dpb_inst_0.INIT_RAM_17 = 256'h4006510E54E5657004839E0439004900EB1522C02F00E254E5C0335200491705;
defparam dpb_inst_0.INIT_RAM_18 = 256'hE1404E50EC5383570E5445B39400E541C57043900EE1B00B257651CDE5445B39;
defparam dpb_inst_0.INIT_RAM_19 = 256'h50E5459C8330049525205839525205C59605A00E54257005441C04356059400E;
defparam dpb_inst_0.INIT_RAM_1A = 256'hC005254E105E950254F0E542143055E00C25C8560142540E5421430455E2504E;
defparam dpb_inst_0.INIT_RAM_1B = 256'h0083530D543930D90E5421705449200429700254F00E5B3A240E5A45E5205441;
defparam dpb_inst_0.INIT_RAM_1C = 256'h4034E5D753005C215721830EFE005DC4393000349E57C03E14000540504E5321;
defparam dpb_inst_0.INIT_RAM_1D = 256'h05C05F3D055139405245105E50A539C94505F00BE12600349E5085522D5E00F2;
defparam dpb_inst_0.INIT_RAM_1E = 256'h5522500C32300A591335320450349E5740542F00A5D25600542200EFE00254D0;
defparam dpb_inst_0.INIT_RAM_1F = 256'h95001045000540A57E18300537218300DF205400571D97C00C25832583054002;
defparam dpb_inst_0.INIT_RAM_20 = 256'h0A00254E594100A5CC9556005404E5D5721830255E94EF3025F0005F002530A5;
defparam dpb_inst_0.INIT_RAM_21 = 256'hB807B84A06062387B042387B82AB07B0B2387B80A0D220EC0F4F6C8E681AA8F8;
defparam dpb_inst_0.INIT_RAM_22 = 256'h6D501E89FAD9709A4018B092A48FB4507B4A0FB6680AA8468F68780A44052387;
defparam dpb_inst_0.INIT_RAM_23 = 256'h92DF3A06284E668197A361F055018BE07BFB001865C3BD3AE3F105E9BBB39469;
defparam dpb_inst_0.INIT_RAM_24 = 256'hFBF07B869CD9FC2D0819DDB092DF30EB3AE30EE81B9CD1B892DF30E0EC0CE830;
defparam dpb_inst_0.INIT_RAM_25 = 256'h5E8239431EA8D030E97B687BA0FBFB913CE130E13F9F9B9947FB1896507BC6B0;
defparam dpb_inst_0.INIT_RAM_26 = 256'hD03FE8060B7743AA8D030E2636702E97A76286E468866E69201EF67A4D03CE00;
defparam dpb_inst_0.INIT_RAM_27 = 256'h9F108B46708B86D00BC6300BB688962F8CE850867A4D03CE33B9E088561E0BAD;
defparam dpb_inst_0.INIT_RAM_28 = 256'h4306A2D48AC27A92FB0B43AADD430E033E980643A2309B2B26682E2B6E1670CA;
defparam dpb_inst_0.INIT_RAM_29 = 256'h0CBD0E1E00707A58F0FB87B0BADD91E0265380655D08A6D870B43F1DAE3CA02D;
defparam dpb_inst_0.INIT_RAM_2A = 256'hE063DAE0CBDF0070CA0C290328F0D266DC40D31A361E06900EEE58730A801EB7;
defparam dpb_inst_0.INIT_RAM_2B = 256'h10B6D86081905115D287B60FB0ED301D97AE304E880ECBDCD0DA0E22E0F2C181;
defparam dpb_inst_0.INIT_RAM_2C = 256'hD00115D021680E2C0EA700E487D1D590014870CA900115D58B6D0313690D115D;
defparam dpb_inst_0.INIT_RAM_2D = 256'h160B8C807B559707F0707F8A037070BDD7DD0708C0077798DB8D070E061D2EE0;
defparam dpb_inst_0.INIT_RAM_2E = 256'h670ED3D3D58F02A0E2CFF022C02A8080EA4628D0FA2650B7D407E0019113AF30;
defparam dpb_inst_0.INIT_RAM_2F = 256'h0330E285EA9F002C2D03A701E0CA7F6B0E2C2D03A777706F1ED0228972E40EEE;
defparam dpb_inst_0.INIT_RAM_30 = 256'hFE0710A2C417CC1001A0068BFC417A34E0524E1131E9F1EC6301F9D01F878F95;
defparam dpb_inst_0.INIT_RAM_31 = 256'hC124190FE407BBC0DC41FC01CEDF6E70E05E207A678B016E70985E407A683937;
defparam dpb_inst_0.INIT_RAM_32 = 256'h16283B387EA806AB9BB086A8FBABCF371C0D571FC81526DCEDFFF910FC0D1754;
defparam dpb_inst_0.INIT_RAM_33 = 256'h43FC38EC01DFE1FF085D5734FF08C4140000FF504400054120451204E5F69082;
defparam dpb_inst_0.INIT_RAM_34 = 256'hF21D43DD1D901E80A29D001FC129DC01E3129DC01E219D0D33F1B22C010ED41D;
defparam dpb_inst_0.INIT_RAM_35 = 256'hFA1F0093BEA2D71DBE5EFF10010D325EFF1D400129DC01F6129D341F2129DC01;
defparam dpb_inst_0.INIT_RAM_36 = 256'hFFFF30B229DC01FE1206DA2093BEA2D51DBEAEFF10010D32AEFF1D400129DC01;
defparam dpb_inst_0.INIT_RAM_37 = 256'hB3C0DE1DBECDAFF1001430E4036A6009B37CDAFF1001770E706F6A3770E706F6;
defparam dpb_inst_0.INIT_RAM_38 = 256'hFD27D70E706F6C17D70E706F6FFFFC99DF01001D409D0019D00198DF3704F009;
defparam dpb_inst_0.INIT_RAM_39 = 256'hF6FFFFBB7D70E706F67DA7D70E706F6FFFF7DE47D70E706F6D37D70E706F6FFF;
defparam dpb_inst_0.INIT_RAM_3A = 256'h0E706F6FFFFA87D70E706F67D77D70E706F6FFFF7D827D70E706F6B17D70E706;
defparam dpb_inst_0.INIT_RAM_3B = 256'h5204E10E97520F40E254E5C033520043540D12039D1E949D17D70E706F6A07D7;
defparam dpb_inst_0.INIT_RAM_3C = 256'h9245200335244104591C03940520CC97045435454032F22509E1049850F40453;
defparam dpb_inst_0.INIT_RAM_3D = 256'h4033524410459694FD081108550390E254410043540B31D00E54492700415200;
defparam dpb_inst_0.INIT_RAM_3E = 256'hA8F9D9F2D0410010EE4B535E0030F8D103F1D138EB31430B31DC9C8804C00435;
defparam dpb_inst_0.INIT_RAM_3F = 256'hE02F3094E140C389109380000000999E1C54FD904DA6FA1431E0F8D163112707;

DPB dpb_inst_1 (
    .DOA({dpb_inst_1_douta_w[11:0],douta[7:4]}),
    .DOB({dpb_inst_1_doutb_w[11:0],doutb[7:4]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7:4]})
);

defparam dpb_inst_1.READ_MODE0 = 1'b0;
defparam dpb_inst_1.READ_MODE1 = 1'b0;
defparam dpb_inst_1.WRITE_MODE0 = 2'b00;
defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
defparam dpb_inst_1.BIT_WIDTH_0 = 4;
defparam dpb_inst_1.BIT_WIDTH_1 = 4;
defparam dpb_inst_1.BLK_SEL_0 = 3'b000;
defparam dpb_inst_1.BLK_SEL_1 = 3'b000;
defparam dpb_inst_1.RESET_MODE = "SYNC";
defparam dpb_inst_1.INIT_RAM_00 = 256'hDA00C41C0003C40C0004C40C0007C40C0005C40C0004C40C000BC40C0315444F;
defparam dpb_inst_1.INIT_RAM_01 = 256'h07666040C9DA2224444404C41C44451804A3F160C7F2021170040100200ED53E;
defparam dpb_inst_1.INIT_RAM_02 = 256'h000000000000000027426667765244527664C9D30029DA000332764233223323;
defparam dpb_inst_1.INIT_RAM_03 = 256'h01015503452BE03006241100C8D0300C8D830FC7C323F128D4E70B200FDD35E0;
defparam dpb_inst_1.INIT_RAM_04 = 256'h001028F328F1102B0CC028F010CC028F45342FC0330020F46302C0003FF7F0BE;
defparam dpb_inst_1.INIT_RAM_05 = 256'h220EC02B4630CCB09C01CBBDBD45342CD5A662715010728A101C8F11D082D092;
defparam dpb_inst_1.INIT_RAM_06 = 256'h42CED138DAF20E343D04202B46342245303B2FE00CEF07CD0920018D031200BC;
defparam dpb_inst_1.INIT_RAM_07 = 256'hEE1A43CF1222CBC300302C03C201C34537CC4020014530003CB4630103CC0003;
defparam dpb_inst_1.INIT_RAM_08 = 256'h2CABE01017553028D03120ECF1212BC3F040202B463CBE15570F030223C3125E;
defparam dpb_inst_1.INIT_RAM_09 = 256'h60402000D0B08E1DE1EC023C3702360060044252502F1121CB753F7CBD2B7020;
defparam dpb_inst_1.INIT_RAM_0A = 256'hF000F0F0EFF000700000D0C08FF0E000F0E0C0CFF0E0D0D0C0B03030F0D0B090;
defparam dpb_inst_1.INIT_RAM_0B = 256'h301020D0C08FF050105010E010C0CFF01000CFF0100000E0F08FF0F0E0F0E0CF;
defparam dpb_inst_1.INIT_RAM_0C = 256'h408FF060E0F0CFF050F0E03030BFF0808070408FF060E040CFF050F0E030BFF0;
defparam dpb_inst_1.INIT_RAM_0D = 256'hF0CFF000F0E03030BFF01000008070408FF0F0E040CFF000F0E030BFF0807070;
defparam dpb_inst_1.INIT_RAM_0E = 256'hCFF030906080807FF0908FF070F0CFF050E030B05FF01000007070408FF0F0E0;
defparam dpb_inst_1.INIT_RAM_0F = 256'h303000C0BFF050A0C0B08FF0A090F0CFF0309060808FF050A0B0B08FF0A09070;
defparam dpb_inst_1.INIT_RAM_10 = 256'h80EFF0807FF0807070401020D0C08FF060E00FF0F0105010E010C0CFF050F0E0;
defparam dpb_inst_1.INIT_RAM_11 = 256'h70E010E0D0D08FF0C0D0D00FF0C0201010C0CFF040D0C04FF0A010A0C0B00FF0;
defparam dpb_inst_1.INIT_RAM_12 = 256'h666402665FF02010D0D0108FF0E01010D0C0CFF0B010C0BFF000D000C0CFF0F0;
defparam dpb_inst_1.INIT_RAM_13 = 256'h2764274027664027666740302676742642667640276427650266664244502666;
defparam dpb_inst_1.INIT_RAM_14 = 256'h7642676402777664077667742766426650222666664264272664026666666740;
defparam dpb_inst_1.INIT_RAM_15 = 256'h4540267642776402666642775266427664026766402766652674276526665026;
defparam dpb_inst_1.INIT_RAM_16 = 256'h7666502664276764266767506664276402766766426752740220767742666502;
defparam dpb_inst_1.INIT_RAM_17 = 256'h4026742666676640276664277402440236667432740237676432776750766526;
defparam dpb_inst_1.INIT_RAM_18 = 256'h6642665266676665266776676402666666427740266640267676764266776676;
defparam dpb_inst_1.INIT_RAM_19 = 256'h5266066666502766764066666764266665275026667650267766777642664026;
defparam dpb_inst_1.INIT_RAM_1A = 256'h6526766642666427664266776752764022766664066774066776752776674266;
defparam dpb_inst_1.INIT_RAM_1B = 256'h0266750667775264066776526776402676502766402666607406677766426776;
defparam dpb_inst_1.INIT_RAM_1C = 256'h5277666665026666667664266402660777503207665262766420274260766764;
defparam dpb_inst_1.INIT_RAM_1D = 256'h2667765206777642677742665276766675274026667402076650776766742767;
defparam dpb_inst_1.INIT_RAM_1E = 256'h7677402245402767677605274207665262677652766764026717526640277420;
defparam dpb_inst_1.INIT_RAM_1F = 256'h7777427420264276666640260676640244527402666642602276667664264027;
defparam dpb_inst_1.INIT_RAM_20 = 256'h4302767666765276666765026427666667664076766766427765027402775276;
defparam dpb_inst_1.INIT_RAM_21 = 256'hC227C30381463026C463027C303424C453025C343413843F301F102FE303F303;
defparam dpb_inst_1.INIT_RAM_22 = 256'h5C020F706C3CB45392B704537025C1025C1024C81313F1113002B38311463024;
defparam dpb_inst_1.INIT_RAM_23 = 256'h06CCD771020F117CCB701CE21F2B70027CCD00001CCD7CD7CDA2203BCDCD7000;
defparam dpb_inst_1.INIT_RAM_24 = 256'h6CA27C0104CCA1BE0C002C0206CCD23CD7CD23126C04C51206CCD0123220F732;
defparam dpb_inst_1.INIT_RAM_25 = 256'h0F7FD7FD8305CFDD3C4CF26CF27CCDCCD03CD13CDAC4CD05C44CA101A26C01A2;
defparam dpb_inst_1.INIT_RAM_26 = 256'hCFDA022EFD50FD705CFDD30100223FCB701020F0102019E7528FDE406CFD0323;
defparam dpb_inst_1.INIT_RAM_27 = 256'hCAA27C01A25C01A26C01B25C0101014120F7029E506CFD13FD7CD1F20E0EFD05;
defparam dpb_inst_1.INIT_RAM_28 = 256'hFD4F7AE1102D003C4CFDFD705CED83FDF07500FD7FD8DCEC1D031FFD80814453;
defparam dpb_inst_1.INIT_RAM_29 = 256'h200C010362B463F14C7CC4CFD05CCCF110C0100C4E9105C44FDEDAEF03C1F2AE;
defparam dpb_inst_1.INIT_RAM_2A = 256'h32E4C31200CA12B453453746375453000702740200002E7C03FF02B403020F75;
defparam dpb_inst_1.INIT_RAM_2B = 256'h120FC004111001EED226C227C07D402DCB03020F020300C75452453034533020;
defparam dpb_inst_1.INIT_RAM_2C = 256'hE030EED4A1914533453B2FF02B7EDE101102B4531021EED220FC061001001EED;
defparam dpb_inst_1.INIT_RAM_2D = 256'h10208C02B7ECC6CE6CECED1F127CEC06C433CEF1F1CE4E123023CE014B2D1F3B;
defparam dpb_inst_1.INIT_RAM_2E = 256'hE407D2D2D51546345334A463346302B45320023453103C0BC02B7462CCE11A40;
defparam dpb_inst_1.INIT_RAM_2F = 256'h121CB022F1CA46300C463480E45341E745300C4634000EE507D4637CB0302FFF;
defparam dpb_inst_1.INIT_RAM_30 = 256'hF34524020A2D0D2001F22EEDD0D2BED634530305C03CC03004024CF18ACB74CF;
defparam dpb_inst_1.INIT_RAM_31 = 256'hB2041F2FF12EED0BC0C2D0E20BC0E7F1D25FE2E00E1E31D7F1025F02E00EDED7;
defparam dpb_inst_1.INIT_RAM_32 = 256'h4CF12EDCB7F24EEDCEDC3EF27CED01CFC0BC082D0E2C00C0BC000E02E0BCEDE0;
defparam dpb_inst_1.INIT_RAM_33 = 256'h8DAED03382F3F3FF4608080CFF460C080222FF050D002676526764266764C463;
defparam dpb_inst_1.INIT_RAM_34 = 256'h03200C032DF20F34304C0C100204C3410E204C3010D2EDBE10F066130123012D;
defparam dpb_inst_1.INIT_RAM_35 = 256'h062E2B72000C072DB553BF0402BE1153BF05540204C34105204C0F109204C381;
defparam dpb_inst_1.INIT_RAM_36 = 256'h1111256604C34106240109CB72000C0A2DB5A3BF0402BE11A3BF05540204C351;
defparam dpb_inst_1.INIT_RAM_37 = 256'h02020F2DB5AA7BF0402FD43020E7F2B7027AA7BF0402724C29C0E72724C29C0E;
defparam dpb_inst_1.INIT_RAM_38 = 256'h1707F24C29C0E707F24C29C0E11117D0F3C0002F030FC400F040D004CA21E2B7;
defparam dpb_inst_1.INIT_RAM_39 = 256'h0E1111707F24C29C0E5E07F24C29C0E11114E707F24C29C0E707F24C29C0E111;
defparam dpb_inst_1.INIT_RAM_3A = 256'h4C29C0E1111717F24C29C0E5E17F24C29C0E11114E017F24C29C0E717F24C29C;
defparam dpb_inst_1.INIT_RAM_3B = 256'h4526642666642652376764327767507765244526666674ED27F24C29C0E727F2;
defparam dpb_inst_1.INIT_RAM_3C = 256'h7776522776766406676677642642666526676676427767742764076742652545;
defparam dpb_inst_1.INIT_RAM_3D = 256'h5277676642666666640644063327426767765277650676422667767522666522;
defparam dpb_inst_1.INIT_RAM_3E = 256'h3C0CCCABE0C0502CFFCDCD0350CC0AC0CC0ACCD1366675067662266226622776;
defparam dpb_inst_1.INIT_RAM_3F = 256'h27764276665223333226200000004442444444C50C000D18D03C0AC08C05CB46;

endmodule //blk_mem_gen_0
