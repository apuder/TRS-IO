//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.9 Beta-4 Education
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Fri Jan 26 20:34:30 2024

module blk_mem_gen_6 (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [7:0] douta;
output [7:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [14:0] ada;
input [7:0] dina;
input [14:0] adb;
input [7:0] dinb;

wire [14:0] dpb_inst_0_douta_w;
wire [0:0] dpb_inst_0_douta;
wire [14:0] dpb_inst_0_doutb_w;
wire [0:0] dpb_inst_0_doutb;
wire [14:0] dpb_inst_1_douta_w;
wire [1:1] dpb_inst_1_douta;
wire [14:0] dpb_inst_1_doutb_w;
wire [1:1] dpb_inst_1_doutb;
wire [14:0] dpb_inst_2_douta_w;
wire [2:2] dpb_inst_2_douta;
wire [14:0] dpb_inst_2_doutb_w;
wire [2:2] dpb_inst_2_doutb;
wire [14:0] dpb_inst_3_douta_w;
wire [3:3] dpb_inst_3_douta;
wire [14:0] dpb_inst_3_doutb_w;
wire [3:3] dpb_inst_3_doutb;
wire [11:0] dpb_inst_4_douta_w;
wire [3:0] dpb_inst_4_douta;
wire [11:0] dpb_inst_4_doutb_w;
wire [3:0] dpb_inst_4_doutb;
wire [14:0] dpb_inst_5_douta_w;
wire [4:4] dpb_inst_5_douta;
wire [14:0] dpb_inst_5_doutb_w;
wire [4:4] dpb_inst_5_doutb;
wire [14:0] dpb_inst_6_douta_w;
wire [5:5] dpb_inst_6_douta;
wire [14:0] dpb_inst_6_doutb_w;
wire [5:5] dpb_inst_6_doutb;
wire [14:0] dpb_inst_7_douta_w;
wire [6:6] dpb_inst_7_douta;
wire [14:0] dpb_inst_7_doutb_w;
wire [6:6] dpb_inst_7_doutb;
wire [14:0] dpb_inst_8_douta_w;
wire [7:7] dpb_inst_8_douta;
wire [14:0] dpb_inst_8_doutb_w;
wire [7:7] dpb_inst_8_doutb;
wire [11:0] dpb_inst_9_douta_w;
wire [7:4] dpb_inst_9_douta;
wire [11:0] dpb_inst_9_doutb_w;
wire [7:4] dpb_inst_9_doutb;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire cea_w;
wire ceb_w;
wire gw_gnd;

assign cea_w = ~wrea & cea;
assign ceb_w = ~wreb & ceb;
assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[14:0],dpb_inst_0_douta[0]}),
    .DOB({dpb_inst_0_doutb_w[14:0],dpb_inst_0_doutb[0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[0]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b1;
defparam dpb_inst_0.READ_MODE1 = 1'b1;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 1;
defparam dpb_inst_0.BIT_WIDTH_1 = 1;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFD0BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFC4BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFC93FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFC97F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFF948FF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_06 = 256'h0000FFFFFFFFFFFE03F17F4FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_07 = 256'h0000FFFFFFFFFFFC00F2FE57FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_08 = 256'h0000FFFFFFFFFFFC08F5FE59FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_09 = 256'h0000FFFFFFFFFFFE09E4FE207FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0A = 256'h0000FFFFFFFFFFFC0AE5FE603FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0B = 256'h0000FFFFFFFFFFFC13E5FE401FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0C = 256'h0000FFFFFFFFFFFC09EBFE0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0D = 256'h0000FFFFFFFFFFF80AE5FC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0E = 256'h0000FFFFFFFFFFF80B47FC0000FE087FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0F = 256'h0000FFFFFFFFFFF805C7FC0000FCAB52451515FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_10 = 256'h0000FFFFFFFFFFF027C7FC0008F910000005AF4D52D28FFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_11 = 256'h0000FFFFFFFFFFF01797F800007D40000000000000005F5F0D72BFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_12 = 256'h0000FFFFFFFFFFE00DAFF81000F1A000000000000000000000002FFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_13 = 256'h0000FFFFFFFFFFF02DAFF8000070A0800000000000000000000017FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_14 = 256'h0000FFFFFFFFFFE0279BF40000FAA0000000000000000000000017FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_15 = 256'h0000FFFFFFFFFFC09B9BF00000F520000290000000000000000017FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_16 = 256'h0000FFFFFFFFFFE08F9FF82001E080000301806300000000000016FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_17 = 256'h0000FFFFFFFFFFC05F5FE80001F20000438180C7008A4000000015FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_18 = 256'h0000FFFFFFFFFF81BB5FE00001F2800043118EE61521110210000EFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_19 = 256'h0000FFFFFFFFFFC1BF3FE04001F540042830AE6000AA10A800000DFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_1A = 256'h0000FFFFFFFFFF811EDFE80001ED500400B886474F894A9500000DFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_1B = 256'h0000FFFFFFFFFF033EFFC60005D0C0100033AEE51FF7FFFFE0080D7FFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_1C = 256'h0000FFFFFFFFFF033DBFC00003E8400021398CE71FF62A8546800EBFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_1D = 256'h0000FFFFFFFFFF027D7FD40007E2000000318EE6AFF6A44556280EBFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_1E = 256'h0000FFFFFFFFFF007DFFDC0C47EA40000009846E0FF6AAEEA6020EBFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_1F = 256'h0000FFFFFFFFFE00BAFFFC0E03F48000003106274FFEA21D56800BBFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_20 = 256'h0000FFFFFFFFFD047BFFB80C07E880000031D4E64FF6A2151680077FFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_21 = 256'h0000FFFFFFFFFE017B7F824C07E88000001094800FF60154268007BFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_22 = 256'h0000FFFFFFFFFC00F3FF650007D4A00000118C070FF60028560007FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_23 = 256'h0000FFFFFFFFFC0AF5FF690007DA2000003084250FFFFFEA1E0007FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_24 = 256'h0000FFFFFFFFF80575FF508097D420000001CCE1090000A84000057FFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_25 = 256'h0000FFFFFFFFF80BF7FF500007DC8000000180A004010400200007FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_26 = 256'h0000FFFFFFFFF803EBFFD0047FD1A00000000070404108200000057FFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_27 = 256'h0000FFFFFFFFF813EBFE9006FF9AA0000000000000000000000007FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_28 = 256'h0000FFFFFFFFF017DBFEB000FF9708000000000000800808000002BFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_29 = 256'h0000FFFFFFFFE825D7FFA2C01FC82A3B0000000000000000000003DFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_2A = 256'h0000FFFFFFFFF007D7FD6F820FDA2A31B50A3F555FA000000000037FFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_2B = 256'h0000FFFFFFFFF00FB7FD4C001FD80000000011D5557B7DBEB57FFF7FFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_2C = 256'h0000FFFFFFFF8097BFFE4A021F5C000000000D0A42ED4000FFFEBBFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_2D = 256'h0000FFFFFFFF00CFBFFA6B003FDC000000000D7E12EE8000000003FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_2E = 256'h0000FFFFFFFF80B73FF9FCC01ED0000000000C7612EDC000000003FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_2F = 256'h0000FFFFFFFFE09433FCF750FF54000000000D2312F74000000001FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_30 = 256'h0000FFFFFFFFE03FBBFE5DD1FF54000010000DAA12F68000000001AFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_31 = 256'h0000FFFFFFFFF05FDF7FD393FF50000000000C667FBF4000000001AFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_32 = 256'h0000FFFFFFFFF83FFFFFE3A3FEA8000000000BD267A4400000000157FFFFFFFF;
defparam dpb_inst_0.INIT_RAM_33 = 256'h0000FFFFFFFFF80FEFFFF853FE68000000000AC26EEDC000000001EFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_34 = 256'h0000FFFFFFFFFC17F7FFFE07FE68000000000AD27F6E8000000001EFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_35 = 256'h0000FFFFFFFFFE0BFFFFFF97FE68000000000B6203B54000000001CFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_36 = 256'h0000FFFFFFFFFE01FBFFFFE7FE68000000000A7C8356C000000000AFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_37 = 256'h0000FFFFFFFFFF01EDFFFFF7FD68000000000B3A0B56C000000000AFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_38 = 256'h0000FFFFFFFFFF80FEFFFFFFFD7000000000197A0BD74000000000AFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_39 = 256'h0000FFFFFFFFFFC0FEFFFFFFFFF8000000001FDE0356C000000000AFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_3A = 256'h0000FFFFFFFFFFE07F7FFFFFFBD8A51F55FA7DAA7F5EC000000000AFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_3B = 256'h0000FFFFFFFFFFF07FBFFFFFFB48F61756AD1D516EFE55F0000000EFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_3C = 256'h0000FFFFFFFFFFF81FFFFFFFFFFFFFFFFFFFFE8AACAEF5FBFF7DFBFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_3D = 256'h0000FFFFFFFFFFF80FDFFFFFFFFFFFFFFFFFFFFFFFFEFBBFF55577FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_3E = 256'h0000FFFFFFFFFFFC07EFFFFFFFFFFFFFFFFFFFFFFF6FFFEEFF7D57FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_3F = 256'h0000FFFFFFFFFFFE07F7FFFFFFFFFFFFFFFFFFFFFFDDF7F7FFFBAFFFFFFFFFFF;

DPB dpb_inst_1 (
    .DOA({dpb_inst_1_douta_w[14:0],dpb_inst_1_douta[1]}),
    .DOB({dpb_inst_1_doutb_w[14:0],dpb_inst_1_doutb[1]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[1]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[1]})
);

defparam dpb_inst_1.READ_MODE0 = 1'b1;
defparam dpb_inst_1.READ_MODE1 = 1'b1;
defparam dpb_inst_1.WRITE_MODE0 = 2'b00;
defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
defparam dpb_inst_1.BIT_WIDTH_0 = 1;
defparam dpb_inst_1.BIT_WIDTH_1 = 1;
defparam dpb_inst_1.BLK_SEL_0 = 3'b000;
defparam dpb_inst_1.BLK_SEL_1 = 3'b000;
defparam dpb_inst_1.RESET_MODE = "SYNC";
defparam dpb_inst_1.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFC03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFE97FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFF07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFF2FF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFF2FF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_06 = 256'h0000FFFFFFFFFFFE044AFE4FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_07 = 256'h0000FFFFFFFFFFFC05A57E27FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_08 = 256'h0000FFFFFFFFFFFC0551FEA1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_09 = 256'h0000FFFFFFFFFFFC01F3FEA0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0A = 256'h0000FFFFFFFFFFFE09737E803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0B = 256'h0000FFFFFFFFFFFC196BFEA01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0C = 256'h0000FFFFFFFFFFF8136AFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0D = 256'h0000FFFFFFFFFFFC13ABFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0E = 256'h0000FFFFFFFFFFF813CAFC0801FD27FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0F = 256'h0000FFFFFFFFFFF837DAFC0000FB5405A8CA5FFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_10 = 256'h0000FFFFFFFFFFF013DBFC00087E5000009240B2AD097FFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_11 = 256'h0000FFFFFFFFFFF02BDBF80000F82000000000000015B0A0F28FFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_12 = 256'h0000FFFFFFFFFFF067B7F80008FC41000000000000000000000037FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_13 = 256'h0000FFFFFFFFFFE047AFF80000FD0000000000000000000000001DFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_14 = 256'h0000FFFFFFFFFFE08F2FF40000F50000000000000000000000001BFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_15 = 256'h0000FFFFFFFFFFE00F6FF00000F84000000000000000000000001BFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_16 = 256'h0000FFFFFFFFFFC05F77F02001FD2000038082630000000000001DFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_17 = 256'h0000FFFFFFFFFFC097BFE80001F52000030180E72220024000000BFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_18 = 256'h0000FFFFFFFFFFC00FBFE00001E9402207319E66404A44A800000B7FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_19 = 256'h0000FFFFFFFFFF801EFFE00001E0000081298AF55551450220000BFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_1A = 256'h0000FFFFFFFFFF80BEBFE80001E08000102094E62A04A54024000BBFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_1B = 256'h0000FFFFFFFFFF806EBFF80005EA000042319EEF4FF7FFFE8A800BFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_1C = 256'h0000FFFFFFFFFF007C7FD40001E540080439AEF74FF68528BE200BFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_1D = 256'h0000FFFFFFFFFF005DBFD40007D54004803198EE0FF611100E800BFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_1E = 256'h0000FFFFFFFFFE02DD3FD40047D480020039D166AFF611D40E800BFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_1F = 256'h0000FFFFFFFFFF027B7F840E03C120000030188F2FF6082C26200EFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_20 = 256'h0000FFFFFFFFFE01FABF800407D280000030C4C80FF608484E200DFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_21 = 256'h0000FFFFFFFFFC0AFAFFBA3C07D4A00000308C404FF6AA028E0007FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_22 = 256'h0000FFFFFFFFFC097EFF990487C98000003904044FF6AA81062005FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_23 = 256'h0000FFFFFFFFFC01777F950007C4800000288C271FFFFA005E10057FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_24 = 256'h0000FFFFFFFFFC11F7FF53008FA9800000018C6500400A01290007FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_25 = 256'h0000FFFFFFFFF811EDFF400007A3400000018060000800810000055FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_26 = 256'h0000FFFFFFFFF812EFFE30007F840000000000E000000104400007FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_27 = 256'h0000FFFFFFFFF025EFFEE000FFA110000000000004022100000006BFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_28 = 256'h0000FFFFFFFFF023EFFEC000FFA0A0000000000000000100900007EFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_29 = 256'h0000FFFFFFFFF007DFFC4F401F33D5E000000000000000000000037FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_2A = 256'h0000FFFFFFFFE02FDFFD4F802F25D5CE5AF7E4ABF0000000000003FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_2B = 256'h0000FFFFFFFFE027DFFD56003F24000000006F2FFFEED7EBDFFF07EFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_2C = 256'h0000FFFFFFFF804FA7FD88023F42000000000AFE03B7E01FFAD5FDDFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_2D = 256'h0000FFFFFFFF0017AFFB92003F20000000000A9513BB8000000002B7FFFFFFFF;
defparam dpb_inst_1.INIT_RAM_2E = 256'h0000FFFFFFFF000F2FFA1D401F2C000000000B9A13B7000000000357FFFFFFFF;
defparam dpb_inst_1.INIT_RAM_2F = 256'h0000FFFFFFFFC02C4FF91E007EA8000000000BFC13AA8000000003BFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_30 = 256'h0000FFFFFFFFE0BEBEFF2C13FEA4000000000AD65BADC000000001FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_31 = 256'h0000FFFFFFFFE05DDFFF8C05FEA8000000000BBE7F55C000000001FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_32 = 256'h0000FFFFFFFFF00F5FBFE403FEA0000000000A3C6EFB8000000001FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_33 = 256'h0000FFFFFFFFF80FEFFFFA83FF90000000000A3E7FBB4000000001BFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_34 = 256'h0000FFFFFFFFFA17F7FFFC53FD90000000000D2C7FDB40000000015FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_35 = 256'h0000FFFFFFFFFC0BF7FFFF87FD98000000000CBC02DFC0000000017FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_36 = 256'h0000FFFFFFFFFF07FBFFFFC7FD80000000000D9603EDC0000000017FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_37 = 256'h0000FFFFFFFFFF81FDFFFFF7FD88000000001CD60BFDC000020000FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_38 = 256'h0000FFFFFFFFFF80FDFFFFFFFE800000000016D6836AC000000000FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_39 = 256'h0000FFFFFFFFFFC17EFFFFFFFD080000400014A2A3FDC000000000FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3A = 256'h0000FFFFFFFFFFE0BF7FFFFFFC275AE0BE80127642B54000000000FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3B = 256'h0000FFFFFFFFFFE02F7FFFFFFCBF4BE8A976F7BED555BE00000000BFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3C = 256'h0000FFFFFFFFFFF03FBFFFFFFFFFFFFFFFB4A177FBFBAAAE55D7556FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3D = 256'h0000FFFFFFFFFFF81FDFFFFFFFFFFFFFFFFFFFFFFB6FDFF6BFFFCBFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3E = 256'h0000FFFFFFFFFFFC0FEFFFFFFFFFFFFFFFFFFFFFEFFEDABBABD7FFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3F = 256'h0000FFFFFFFFFFFE07E7FFFFFFFFFFFFFFFFFFFFFFF7BDDDAAAEFFFFFFFFFFFF;

DPB dpb_inst_2 (
    .DOA({dpb_inst_2_douta_w[14:0],dpb_inst_2_douta[2]}),
    .DOB({dpb_inst_2_doutb_w[14:0],dpb_inst_2_doutb[2]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[2]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[2]})
);

defparam dpb_inst_2.READ_MODE0 = 1'b1;
defparam dpb_inst_2.READ_MODE1 = 1'b1;
defparam dpb_inst_2.WRITE_MODE0 = 2'b00;
defparam dpb_inst_2.WRITE_MODE1 = 2'b00;
defparam dpb_inst_2.BIT_WIDTH_0 = 1;
defparam dpb_inst_2.BIT_WIDTH_1 = 1;
defparam dpb_inst_2.BLK_SEL_0 = 3'b000;
defparam dpb_inst_2.BLK_SEL_1 = 3'b000;
defparam dpb_inst_2.RESET_MODE = "SYNC";
defparam dpb_inst_2.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFC97FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFD0BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFC57FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFC97FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFDA97F3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_06 = 256'h0000FFFFFFFFFFFFF7F17F1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_07 = 256'h0000FFFFFFFFFFFC0272FE47FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_08 = 256'h0000FFFFFFFFFFFC08F6FE59FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_09 = 256'h0000FFFFFFFFFFFE0955FE20FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0A = 256'h0000FFFFFFFFFFFC05E5FE207FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0B = 256'h0000FFFFFFFFFFFC15C5FC401FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0C = 256'h0000FFFFFFFFFFFC15C3FE0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0D = 256'h0000FFFFFFFFFFF80AEAFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0E = 256'h0000FFFFFFFFFFF805CFFC0803FD5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0F = 256'h0000FFFFFFFFFFF00347FC00007C0AA81221FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_10 = 256'h0000FFFFFFFFFFF825C7FC00007880000A68AB4D5897FFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_11 = 256'h0000FFFFFFFFFFF00587FA0000FAD0000000000002D6CF5F5D7FFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_12 = 256'h0000FFFFFFFFFFF00BCFF80008F29000000000000000000000005FFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_13 = 256'h0000FFFFFFFFFFE05BABF80000F051400000000000000000000017FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_14 = 256'h0000FFFFFFFFFFE04BBFF80000F0A0000000000000000000000017FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_15 = 256'h0000FFFFFFFFFFC0AD9FF00000F500000000000000000000000015FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_16 = 256'h0000FFFFFFFFFFC08F9FF02000F240000299806700000000000013FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_17 = 256'h0000FFFFFFFFFFC09F6FF80001E88001000086470800000000001EFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_18 = 256'h0000FFFFFFFFFF81BE5FE80001F2000042018EE72510120120000DFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_19 = 256'h0000FFFFFFFFFF81B75FE00023F5401010101A0722042A5084000EFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1A = 256'h0000FFFFFFFFFF812EBFE00001EA4000800AAEE550AA102A81000EFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1B = 256'h0000FFFFFFFFFF033CFFC40005E5400200258A070FF7FFC120000EFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1C = 256'h0000FFFFFFFFFF032FBFD40001D2400080399CE51FF668921E000EBFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1D = 256'h0000FFFFFFFFFF037D7FC80003E8400008398686AFF6AAA556200EBFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1E = 256'h0000FFFFFFFFFF007DFFD40003E240000021C0175FF6A5CAB6080EBFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1F = 256'h0000FFFFFFFFFE04FCFFFC0603EA8000000804000FF6A30E8E800BDFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_20 = 256'h0000FFFFFFFFFE067B7FFC0E07E8A00000208CE04FF6A3C2A680077FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_21 = 256'h0000FFFFFFFFFE00BBFFA20407C2800000318CC72FF600502688057FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_22 = 256'h0000FFFFFFFFFC01F3FFA3048FD2000000398C662FF600281680077FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_23 = 256'h0000FFFFFFFFFA0DF5FF610007AAA00000298CD03FF7C0152E0007DFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_24 = 256'h0000FFFFFFFFF80AF57F40008FD4200000110CE6102AA054000006DFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_25 = 256'h0000FFFFFFFFF80AF7FF700007D42000000100E512402010000007FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_26 = 256'h0000FFFFFFFFF40BEBFFD0047FBBA0000000006008082000000006BFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_27 = 256'h0000FFFFFFFFF803EBFE1002FF8D40000000000000000000000005FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_28 = 256'h0000FFFFFFFFF007DBFE3000FF5D10000000000002000020000002BFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_29 = 256'h0000FFFFFFFFF033D7FFA1C03FC02A000000000000011000000003FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2A = 256'h0000FFFFFFFFF007D7FDAB802FCA2A31A5485BFE80000000000003DFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2B = 256'h0000FFFFFFFFF00F97FD63003FDA0000000FD8F55555AD56FFC0037FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2C = 256'h0000FFFFFFFF800FBFFD54002F58000000000FAA42EAA3FEAF7F5F7FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2D = 256'h0000FFFFFFFF008FBFFA75003F4C000000000DEA42E50000000007FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2E = 256'h0000FFFFFFFF009FBFFBFD405F50000000000D6412EAC000000003FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2F = 256'h0000FFFFFFFFC09F17FCDF407F54000000000C4A1ADDC0000000016FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_30 = 256'h0000FFFFFFFFC0B7BFFE5B89FF54000000000D2A12DB0000000001B7FFFFFFFF;
defparam dpb_inst_2.INIT_RAM_31 = 256'h0000FFFFFFFFE05FBFFF9383FF54000000000C5242EB0000000001B7FFFFFFFF;
defparam dpb_inst_2.INIT_RAM_32 = 256'h0000FFFFFFFFF03FDFFFE333FF58000000000DD67FAEC000000001AFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_33 = 256'h0000FFFFFFFFF80FEFFFF0B3FC68000000000DD47ED680000000016FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_34 = 256'h0000FFFFFFFFFC17F7FFFE87FE68000000000AF66EADC000000001F7FFFFFFFF;
defparam dpb_inst_2.INIT_RAM_35 = 256'h0000FFFFFFFFFE07F7FFFF17FE60000000000BD60368C000000001B7FFFFFFFF;
defparam dpb_inst_2.INIT_RAM_36 = 256'h0000FFFFFFFFFE03FBFFFFE7FE68000000000B6A02BB4000000000D7FFFFFFFF;
defparam dpb_inst_2.INIT_RAM_37 = 256'h0000FFFFFFFFFF01FDFFFFF7FE6800000000076A2B574000000000AFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_38 = 256'h0000FFFFFFFFFF80FDFFFFFFFD70000000000B2A03BDC000000000AFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_39 = 256'h0000FFFFFFFFFFC0EEFFFFFFFD70000040001B7E02AB4000000000AFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3A = 256'h0000FFFFFFFFFFE07F7FFFFFFBD8A51FA0001FAE03EBC000000000AFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3B = 256'h0000FFFFFFFFFFF03FBFFFFFFBC0B41F56A989552BEAE000000000D7FFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3C = 256'h0000FFFFFFFFFFF81DBFFFFFFFFFFFFFD6AB5EA956955F5BAAAAFFDFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3D = 256'h0000FFFFFFFFFFF80F5FFFFFFFFFFFFFFFFFFFFFDFFF76DFEA843DFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3E = 256'h0000FFFFFFFFFFFC0FEFFFFFFFFFFFFFFFFFFFFEFFFFFFFEFD7D57FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3F = 256'h0000FFFFFFFFFFFE07FFFFFFFFFFFFFFFFFFFFFFFDFFEF777FDBB7FFFFFFFFFF;

DPB dpb_inst_3 (
    .DOA({dpb_inst_3_douta_w[14:0],dpb_inst_3_douta[3]}),
    .DOB({dpb_inst_3_doutb_w[14:0],dpb_inst_3_doutb[3]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[3]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[3]})
);

defparam dpb_inst_3.READ_MODE0 = 1'b1;
defparam dpb_inst_3.READ_MODE1 = 1'b1;
defparam dpb_inst_3.WRITE_MODE0 = 2'b00;
defparam dpb_inst_3.WRITE_MODE1 = 2'b00;
defparam dpb_inst_3.BIT_WIDTH_0 = 1;
defparam dpb_inst_3.BIT_WIDTH_1 = 1;
defparam dpb_inst_3.BLK_SEL_0 = 3'b000;
defparam dpb_inst_3.BLK_SEL_1 = 3'b000;
defparam dpb_inst_3.RESET_MODE = "SYNC";
defparam dpb_inst_3.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFE03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFE47FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFF8BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFF52FF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_06 = 256'h0000FFFFFFFFFFFFF8AAFE5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_07 = 256'h0000FFFFFFFFFFFC04E9FEA7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_08 = 256'h0000FFFFFFFFFFFC05B1FEA3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_09 = 256'h0000FFFFFFFFFFFC00F2FEA4FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0A = 256'h0000FFFFFFFFFFFE0AB37E807FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0B = 256'h0000FFFFFFFFFFFC12EB7E801FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0C = 256'h0000FFFFFFFFFFFC12EBFC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0D = 256'h0000FFFFFFFFFFFC13EBFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0E = 256'h0000FFFFFFFFFFF81B6BFC0803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0F = 256'h0000FFFFFFFFFFF835DBFC08007EE556E89FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_10 = 256'h0000FFFFFFFFFFF027DBFC00007F5001A49050B2C87FFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_11 = 256'h0000FFFFFFFFFFF037DBF800007D0000000000002D2930A1A3FFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_12 = 256'h0000FFFFFFFFFFE06697F80008FD200000000000000000000025EBFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_13 = 256'h0000FFFFFFFFFFF026BFF81000FDA000000000000000000000001BFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_14 = 256'h0000FFFFFFFFFFE02FAFF40000FA4000000000000000000000001DFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_15 = 256'h0000FFFFFFFFFFE00F6FF00000F24000000000000000000000001FFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_16 = 256'h0000FFFFFFFFFFE0576FF02002F4800002988C630000000000001EFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_17 = 256'h0000FFFFFFFFFFC04D5FE80000F520000018C4F600902000000005FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_18 = 256'h0000FFFFFFFFFFC00FBFE00003E940000B014E470845405000000AFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_19 = 256'h0000FFFFFFFFFFC01EBFE04003E2800244500004885280AA0000097FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_1A = 256'h0000FFFFFFFFFF813EDFE00001E5104004A18EEF05514A9420000B7FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_1B = 256'h0000FFFFFFFFFF805EBFFC0003D040100803DA275FFFFE2495000B7FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_1C = 256'h0000FFFFFFFFFF007C7FC80001E8400000014E074FF695459E800BFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_1D = 256'h0000FFFFFFFFFF005D7FD40007D2400000280A560FF64408A6800BFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_1E = 256'h0000FFFFFFFFFE015D7FD40003D5000040018E842FF608C106900BFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_1F = 256'h0000FFFFFFFFFE00BB7F840A03D4400008119E68AFF609D826000EFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_20 = 256'h0000FFFFFFFFFE00FAFF800607C68000000188E20FFE085016000DFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_21 = 256'h0000FFFFFFFFFC0AFAFF9A1C0BE8800000118C860FF65505560007FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_22 = 256'h0000FFFFFFFFFC08FAFFAD0C0FC8A000003000F70FF6AA82A60007FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_23 = 256'h0000FFFFFFFFFC02F6FF9D0007D1000000018CA01FF78240060006FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_24 = 256'h0000FFFFFFFFFC11F7FF35008FC1800000310C6005000500140007FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_25 = 256'h0000FFFFFFFFF813F5FF00000F8980000001C04700008200440006BFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_26 = 256'h0000FFFFFFFFF812EFFE20143FC44000000000E041010440000005DFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_27 = 256'h0000FFFFFFFFF015EFFEF000FFA2A0000000006000000000000007BFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_28 = 256'h0000FFFFFFFFF033EFFED000FFA2A8000000000000001004000007FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_29 = 256'h0000FFFFFFFFF00FDBFE57403FA2C00000000000004000000000035FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2A = 256'h0000FFFFFFFFE057DFFC4DC02F35D5CE5AB7AEA0000000000000037FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2B = 256'h0000FFFFFFFFE047DFFD17001F020000017A679AAABB7AFFE80003FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2C = 256'h0000FFFFFFFFC057AFFD54003F2400000000085D7FBF7FEBFBD5F7FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2D = 256'h0000FFFFFFFF0057AFFA95021F70000000000B3E1BBF8000000007BFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2E = 256'h0000FFFFFFFF002F2FFA1D005EA8000000000ABE53BD8000000002AFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2F = 256'h0000FFFFFFFFC02D2FF91A203EA4000000000BB60BB70000000003FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_30 = 256'h0000FFFFFFFFE0BFBFFE2A23FEA4000000000AFE53B6C000000001FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_31 = 256'h0000FFFFFFFFF05FDF7F2C23FEA0000000000BAC43BEC000000001FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_32 = 256'h0000FFFFFFFFF01FDFFFEC03FEA0000000000A2A66DB0000000001FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_33 = 256'h0000FFFFFFFFF80EEFFFFA83FF90000000000A2A6FADC000000001FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_34 = 256'h0000FFFFFFFFF807E7FFFC23FD90000000000B4A67D640000000015FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_35 = 256'h0000FFFFFFFFFC0BF7FFFF07FD98000000000D2C03B740000000015FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_36 = 256'h0000FFFFFFFFFE03DBFFFFC7FD88000010000CBC036EC000000001BFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_37 = 256'h0000FFFFFFFFFF05FBFFFFF7FD8000000000199E0BAAC000000000FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_38 = 256'h0000FFFFFFFFFF80FDFFFFFFFD80000000001DFE03574000000000FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_39 = 256'h0000FFFFFFFFFFA0FEFFFFFFFE800000400016CA8356C000000000FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_3A = 256'h0000FFFFFFFFFFC0FF7FFFFFFE275BE8000014F202BEC000000000FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_3B = 256'h0000FFFFFFFFFFE07F7FFFFFFE3F5BE0ABF67EAEFF5FA000000000FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_3C = 256'h0000FFFFFFFFFFF03FBFFFFFFFFFFFFAA955A9DEBB6EA9F6FF7FFB7FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_3D = 256'h0000FFFFFFFFFFF81FDFFFFFFFFFFFFFFFFFFFFFFFFBFFFBBDFBEAFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_3E = 256'h0000FFFFFFFFFFFC0FEFFFFFFFFFFFFFFFFFFFFFFF6DBF6FAFD7BFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_3F = 256'h0000FFFFFFFFFFFE07EFFFFFFFFFFFFFFFFFFFFFFFBF7FFFF7FFFFFFFFFFFFFF;

DPB dpb_inst_4 (
    .DOA({dpb_inst_4_douta_w[11:0],dpb_inst_4_douta[3:0]}),
    .DOB({dpb_inst_4_doutb_w[11:0],dpb_inst_4_doutb[3:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[14],ada[13],ada[12]}),
    .BLKSELB({adb[14],adb[13],adb[12]}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[3:0]})
);

defparam dpb_inst_4.READ_MODE0 = 1'b1;
defparam dpb_inst_4.READ_MODE1 = 1'b1;
defparam dpb_inst_4.WRITE_MODE0 = 2'b00;
defparam dpb_inst_4.WRITE_MODE1 = 2'b00;
defparam dpb_inst_4.BIT_WIDTH_0 = 4;
defparam dpb_inst_4.BIT_WIDTH_1 = 4;
defparam dpb_inst_4.BLK_SEL_0 = 3'b100;
defparam dpb_inst_4.BLK_SEL_1 = 3'b100;
defparam dpb_inst_4.RESET_MODE = "SYNC";
defparam dpb_inst_4.INIT_RAM_00 = 256'hBFBD7F5F5F5F5FAFAF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFE7FF6FF6F6FDF6FBFAFBFDBF;
defparam dpb_inst_4.INIT_RAM_02 = 256'h000008FFFFFF1EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_03 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5;
defparam dpb_inst_4.INIT_RAM_04 = 256'hBF5FBFBFBFAFAFAFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFBFFEFBFFDFBFDF6F6FBFBFAFBFAF;
defparam dpb_inst_4.INIT_RAM_06 = 256'h500000AFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_07 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_08 = 256'h5F6BEBEBEBEBEBEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFDF7EFBFFBF6FDFBFDFDFA7F5F6F;
defparam dpb_inst_4.INIT_RAM_0A = 256'hF100000FFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_0B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_0C = 256'hD7D7D7D7DFAFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFBFFDFFFBFEFDFFDFBFE7BFEDFAFD7;
defparam dpb_inst_4.INIT_RAM_0E = 256'hFF100006DFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_0F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_10 = 256'h7E7E7D7E7E7EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFDFFEF7FEFDFBFE7FBFBE7F5F6F5E7E;
defparam dpb_inst_4.INIT_RAM_12 = 256'hFFF00000BEFFFFF2EFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_13 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_14 = 256'hD7D7D6FAFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFDF7FBFDF7EBFDFDFBEBF7DF6D7;
defparam dpb_inst_4.INIT_RAM_16 = 256'hFFFB000005FFFFFF0FFFFFFFFFBFFFF7FFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_17 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_18 = 256'hD7D7D7D7EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFDFF7EFF6FBFD7EBEBEBF6F6FAF6D7D7;
defparam dpb_inst_4.INIT_RAM_1A = 256'hFFFF500000AFFFFFF0FFFFFEFFFF7FFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1C = 256'hBFDFFF1F5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFDF7FFBFEFBE7D7DF6F5F6FBF6BEBEF;
defparam dpb_inst_4.INIT_RAM_1E = 256'hFFFFF0000004FFFFF70FFFF7FFBFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_20 = 256'hF6FFABAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFDFFBFFFE7FBFBF6FDF6FDF6F5FBF5FFA;
defparam dpb_inst_4.INIT_RAM_22 = 256'hFFFFFFB000004FFFFF5EFFFFBFE7FFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_23 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_24 = 256'hFFEAEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFF7FFEFFDF7EFD7FF6FDFDF5FDF5FDFD7DF5FDFD;
defparam dpb_inst_4.INIT_RAM_26 = 256'hFFFFFFFF520000FFFFF1EFFDFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_27 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_28 = 256'hCE9B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFEF7DF7DFDFBF6FDFDF5FDF7DFAFAFE7EBF;
defparam dpb_inst_4.INIT_RAM_2A = 256'hFFFFFFFFF520000FFFBF0FFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFE7FDF6F6FDFBF5FD7D7D6FAF6F5F5F5FB;
defparam dpb_inst_4.INIT_RAM_2E = 256'hFFFFFFFFFF50000CF7DFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFDFFBFFEFDFBFEBF7DFDBEFAFAFAFA7F5F5F5F7F;
defparam dpb_inst_4.INIT_RAM_32 = 256'hFFFFFFFFFFF21000CF6FD78FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_33 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFBFFBFEFBFFDF6FBEFDFAFBEBFD7F5FBFBFFFFF;
defparam dpb_inst_4.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFF77DBFFF78FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_37 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFF7BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DPB dpb_inst_5 (
    .DOA({dpb_inst_5_douta_w[14:0],dpb_inst_5_douta[4]}),
    .DOB({dpb_inst_5_doutb_w[14:0],dpb_inst_5_doutb[4]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[4]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[4]})
);

defparam dpb_inst_5.READ_MODE0 = 1'b1;
defparam dpb_inst_5.READ_MODE1 = 1'b1;
defparam dpb_inst_5.WRITE_MODE0 = 2'b00;
defparam dpb_inst_5.WRITE_MODE1 = 2'b00;
defparam dpb_inst_5.BIT_WIDTH_0 = 1;
defparam dpb_inst_5.BIT_WIDTH_1 = 1;
defparam dpb_inst_5.BLK_SEL_0 = 3'b000;
defparam dpb_inst_5.BLK_SEL_1 = 3'b000;
defparam dpb_inst_5.RESET_MODE = "SYNC";
defparam dpb_inst_5.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFE17FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFC8BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFC17FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFCA7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFE87F3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_06 = 256'h0000FFFFFFFFFFFFFB697F1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_07 = 256'h0000FFFFFFFFFFFC02B2FF47FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_08 = 256'h0000FFFFFFFFFFFC00F5BE53FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_09 = 256'h0000FFFFFFFFFFFE0DA5FE4CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0A = 256'h0000FFFFFFFFFFFE09E5FE207FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0B = 256'h0000FFFFFFFFFFFE0965FE601FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0C = 256'h0000FFFFFFFFFFFC05E5FE000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0D = 256'h0000FFFFFFFFFFF80AA5FC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0E = 256'h0000FFFFFFFFFFFC01C5FC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0F = 256'h0000FFFFFFFFFFF803C6FC08007D1801057FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_10 = 256'h0000FFFFFFFFFFF81347FC00007800325B448F4807FFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_11 = 256'h0000FFFFFFFFFFF002D7FC00007A50000000000552D6CF5E5FFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_12 = 256'h0000FFFFFFFFFFF00FDBF81000784100000000000000000003DFBFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_13 = 256'h0000FFFFFFFFFFE04F8FF80000F001000000000000000000000017FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_14 = 256'h0000FFFFFFFFFFE04B2FFC0001F500000000000000000000000017FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_15 = 256'h0000FFFFFFFFFFE0D79BF40000F500000000000000000000000015FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_16 = 256'h0000FFFFFFFFFFC08F9FF00000F520000298886000000000000015FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_17 = 256'h0000FFFFFFFFFFC09FBFF80000F240004299CC222002000000001BFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_18 = 256'h0000FFFFFFFFFFC1BF6FE00002F4A009423990E74110028000001FFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_19 = 256'h0000FFFFFFFFFF81B76FE00001F420000031C01622A82A0020000FFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_1A = 256'h0000FFFFFFFFFF80B6BFE00001E840024019DC60AA04A52108000DFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_1B = 256'h0000FFFFFFFFFF033EBFC40023EA00004111CC4B3FFF408240400DFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_1C = 256'h0000FFFFFFFFFF033FBFD40003E50011110114071FF602A87E000EFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_1D = 256'h0000FFFFFFFFFF027DBFD40003E5400801082CE6AFF691A20E080EBFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_1E = 256'h0000FFFFFFFFFF007DBFC80003E0800400001C568FF6A3D456200EBFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_1F = 256'h0000FFFFFFFFFF047DBFFC060BE18002003188E00FF6A15E96A00D7FFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_20 = 256'h0000FFFFFFFFFE04BBBFFC0E03E90000080180A74FFEA2A54690077FFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_21 = 256'h0000FFFFFFFFFE057B7FA4040FD6A00000119CE64FF6802806A006FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_22 = 256'h0000FFFFFFFFFE01B3FF930407D68000002000065FF6002806A0057FFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_23 = 256'h0000FFFFFFFFFC0975FF61000FE6A00000018CE0AFF7A8A9568007DFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_24 = 256'h0000FFFFFFFFF80AF5FF49000FAA200000308CE000055005FE00055FFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_25 = 256'h0000FFFFFFFFFC09F7FF700007D22000000080E504120802000005FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_26 = 256'h0000FFFFFFFFF803FBFFD0141F9120000000006000200002000007FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_27 = 256'h0000FFFFFFFFF803EAFE9004FFD91000000000E002110000000006EFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_28 = 256'h0000FFFFFFFFF80BEBFEB000FF9508000000000000000200000002BFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_29 = 256'h0000FFFFFFFFF003D7FDA0C07F5D20000000000004080100000003FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_2A = 256'h0000FFFFFFFFF007D7FFA3402FCA2A31AD5AF00000000000000003FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_2B = 256'h0000FFFFFFFFF02FD7FDE7800FD800009EAF9A6FFFEEAFBE000003DFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_2C = 256'h0000FFFFFFFFE00FB7FD54003F5A000000000FB660D5DEBEAD7F7DDFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_2D = 256'h0000FFFFFFFF008FB7FA64021F08000000000CD51AEA800000000DF7FFFFFFFF;
defparam dpb_inst_5.INIT_RAM_2E = 256'h0000FFFFFFFF0097BFFAF9005F54000000000DD41AE74000000003FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_2F = 256'h0000FFFFFFFFC0975FF9FA201F54000000000D6A0AEAC000000002F7FFFFFFFF;
defparam dpb_inst_5.INIT_RAM_30 = 256'h0000FFFFFFFFE0BEBBFCDE89FF54000000000D9412ED8000000001AFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_31 = 256'h0000FFFFFFFFE03BBFFF93ABFF54000000000CF602D58000000001AFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_32 = 256'h0000FFFFFFFFF01DDEFFC38BFE58000000000ADE67B5C0000200016FFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_33 = 256'h0000FFFFFFFFF82FEFFFF123FE68000000000BD666FB4000000001D7FFFFFFFF;
defparam dpb_inst_5.INIT_RAM_34 = 256'h0000FFFFFFFFFC17FFFFFCC7FE68000000000CB66EAB8000000001F7FFFFFFFF;
defparam dpb_inst_5.INIT_RAM_35 = 256'h0000FFFFFFFFFE07F7FFFF27FE60000000000AF642DAC000000001F7FFFFFFFF;
defparam dpb_inst_5.INIT_RAM_36 = 256'h0000FFFFFFFFFE0BFBFFFFC7FE70000030000BD623DB8000000000EFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_37 = 256'h0000FFFFFFFFFF01FDFFFFE7FE68000000000E6A8AFFC000000000AFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_38 = 256'h0000FFFFFFFFFF81FDFFFFFFFE700000000002522AFBC000000000AFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_39 = 256'h0000FFFFFFFFFFC0FEFFFFFFFD70000000001D3603FDC000000000AFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_3A = 256'h0000FFFFFFFFFFE06F7FFFFFFDD8F40000001B4E83D54000000000AFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_3B = 256'h0000FFFFFFFFFFE0377FFFFFF9D0A51F544BD1F5F9B56000000000AFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_3C = 256'h0000FFFFFFFFFFF05FBFFFFFFFFFFE8556EA76B355B5FEAD55FE81D7FFFFFFFF;
defparam dpb_inst_5.INIT_RAM_3D = 256'h0000FFFFFFFFFFF81FDFFFFFFFFFFFFFFFFFFFFFFFFFABA45256D77FFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_3E = 256'h0000FFFFFFFFFFF80FDFFFFFFFFFFFFFFFFFFFFFF7FFEFFBFABAEBFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_3F = 256'h0000FFFFFFFFFFFC07AFFFFFFFFFFFFFFFFFFFFEEFF5F5555D555FFFFFFFFFFF;

DPB dpb_inst_6 (
    .DOA({dpb_inst_6_douta_w[14:0],dpb_inst_6_douta[5]}),
    .DOB({dpb_inst_6_doutb_w[14:0],dpb_inst_6_doutb[5]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[5]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[5]})
);

defparam dpb_inst_6.READ_MODE0 = 1'b1;
defparam dpb_inst_6.READ_MODE1 = 1'b1;
defparam dpb_inst_6.WRITE_MODE0 = 2'b00;
defparam dpb_inst_6.WRITE_MODE1 = 2'b00;
defparam dpb_inst_6.BIT_WIDTH_0 = 1;
defparam dpb_inst_6.BIT_WIDTH_1 = 1;
defparam dpb_inst_6.BLK_SEL_0 = 3'b000;
defparam dpb_inst_6.BLK_SEL_1 = 3'b000;
defparam dpb_inst_6.RESET_MODE = "SYNC";
defparam dpb_inst_6.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFF03FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFF4BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFF1BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFB3FF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_06 = 256'h0000FFFFFFFFFFFFFAF2FF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_07 = 256'h0000FFFFFFFFFFFC04E5FE27FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_08 = 256'h0000FFFFFFFFFFFC0552FEA3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_09 = 256'h0000FFFFFFFFFFFC00F1FEA1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0A = 256'h0000FFFFFFFFFFFC0552FEA07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0B = 256'h0000FFFFFFFFFFFC05D3FE803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0C = 256'h0000FFFFFFFFFFFC196BFD400FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0D = 256'h0000FFFFFFFFFFFC11EBFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0E = 256'h0000FFFFFFFFFFF817EBFC0803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0F = 256'h0000FFFFFFFFFFF836DBFC08007D42AA17FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_10 = 256'h0000FFFFFFFFFFF025DBFC00007EE98CA42950027FFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_11 = 256'h0000FFFFFFFFFFF02FCBF800007D4000000000B2AD2930A9FFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_12 = 256'h0000FFFFFFFFFFF063A7F8000076900000000000000000005D6A57FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_13 = 256'h0000FFFFFFFFFFF057B7FC10017D4000000000000000000000001DFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_14 = 256'h0000FFFFFFFFFFE02FAFF40000F8A000000000000000000000001BFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_15 = 256'h0000FFFFFFFFFFC02F6FF00000F8A000000000000000000000001BFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_16 = 256'h0000FFFFFFFFFFE05B7FF00011F080000108C4000000000000001BFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_17 = 256'h0000FFFFFFFFFFC0575FE82000E8800003914C020200000000000EFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_18 = 256'h0000FFFFFFFFFFA00B9FE00003EA000003180E202A0408020000057FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_19 = 256'h0000FFFFFFFFFFC01EDFE00001E28020502994C74902815500000AFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_1A = 256'h0000FFFFFFFFFF811EBFE00003F280080829ACEF10AA10CAA0800AFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_1B = 256'h0000FFFFFFFFFF8076FFF80003E54004003191609FFC956928000AFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_1C = 256'h0000FFFFFFFFFF806C7FD80003D0400000094E774FF755017E000BBFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_1D = 256'h0000FFFFFFFFFF013D7FC80043D0400080210C804FF72A5556800BFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_1E = 256'h0000FFFFFFFFFF00BD7FD40003D6400000380EEE6FF61482AE400BFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_1F = 256'h0000FFFFFFFFFE02D97F840443CA4000002100AEAFF615CC46000BFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_20 = 256'h0000FFFFFFFFFE02FA7F840E03D4C000003194050FF6094E16000DFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_21 = 256'h0000FFFFFFFFFC00FAFFA80C0BC0000000319C060FF60880A6000DBFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_22 = 256'h0000FFFFFFFFFC08FAFFAC4C07C0800000280C040FF65501560007FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_23 = 256'h0000FFFFFFFFFC05F6FF99000F88000000000C000FF705000610057FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_24 = 256'h0000FFFFFFFFFC05F77F520007D480000031886000F001FFFE4007FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_25 = 256'h0000FFFFFFFFF81375FF400017AD800000000067110020A8100007FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_26 = 256'h0000FFFFFFFFF819EDFE20101FAA8000000000E0220249104000077FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_27 = 256'h0000FFFFFFFFF015EFFEB002FFA4A0000000001020002000000005FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_28 = 256'h0000FFFFFFFFF027EFFEB000FFA968000000000000000000800007EFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_29 = 256'h0000FFFFFFFFF035EFFE5780FFA200000000000000008000000002FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_2A = 256'h0000FFFFFFFFE02BDFFC4DC00F25D5CED2ED0000000001000000035FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_2B = 256'h0000FFFFFFFFE047DFFC17820F0500076BD16DD55555FFC00000037FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_2C = 256'h0000FFFFFFFFE047AFFD50001FA0000000000AED017B75D5FFD5D77FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_2D = 256'h0000FFFFFFFF0017AFFB8A021F74000000000BAA53B500000000BF7FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_2E = 256'h0000FFFFFFFF000F2FFA9A805F28000000000B2E5BBA80000000036FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_2F = 256'h0000FFFFFFFFC02E2FFA1EA01EA4000000000ADC13BD80000000035FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_30 = 256'h0000FFFFFFFFC0B7BEFE3EA1FEA4000000000A6A53B74000000001FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_31 = 256'h0000FFFFFFFFE05FBDFF2C03FEA0000000000B0A03AB4000000001FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_32 = 256'h0000FFFFFFFFE85FDFEFCC03FFA0000000000DAA7EEF0000020001FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_33 = 256'h0000FFFFFFFFF00FEFFFF413FD90000000000C3A6FAEC0000000017FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_34 = 256'h0000FFFFFFFFF807EFFFFC23FD90000000000B5A6FBEC0000000015FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_35 = 256'h0000FFFFFFFFFC0FD7FFFE03FD88000000000D9A7F6FC0000000014FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_36 = 256'h0000FFFFFFFFFE0BFBFFFF87FD88000000000D2A03754000000001BFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_37 = 256'h0000FFFFFFFFFF01FBFFFFE7FD900000000015BE0B554000000000FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_38 = 256'h0000FFFFFFFFFF80FDFFFFFFFD80000000001FAE0BAD4000000000FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_39 = 256'h0000FFFFFFFFFF80FEFFFFFFFD800000000013EA82AB4000000000FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_3A = 256'h0000FFFFFFFFFFC0FEFFFFFFFA270000000016BA82ABC000000000FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_3B = 256'h0000FFFFFFFFFFE07F7FFFFFFE2F5AE0AFBD2F1B00EEC000000000FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_3C = 256'h0000FFFFFFFFFFF03FBFFFFFFFFF097ABB1FCBCDEEEAAB5BBFC000BFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_3D = 256'h0000FFFFFFFFFFF81FDFFFFFFFFFFFFFFFFFFFFFFFFBFC7BEFBD7EBFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_3E = 256'h0000FFFFFFFFFFFC0FFFFFFFFFFFFFFFFFFFFFFFFFF77D5D6FEFBFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_3F = 256'h0000FFFFFFFFFFFE07EFFFFFFFFFFFFFFFFFFFFFFFFFDFFFF7FFF7FFFFFFFFFF;

DPB dpb_inst_7 (
    .DOA({dpb_inst_7_douta_w[14:0],dpb_inst_7_douta[6]}),
    .DOB({dpb_inst_7_doutb_w[14:0],dpb_inst_7_doutb[6]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[6]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[6]})
);

defparam dpb_inst_7.READ_MODE0 = 1'b1;
defparam dpb_inst_7.READ_MODE1 = 1'b1;
defparam dpb_inst_7.WRITE_MODE0 = 2'b00;
defparam dpb_inst_7.WRITE_MODE1 = 2'b00;
defparam dpb_inst_7.BIT_WIDTH_0 = 1;
defparam dpb_inst_7.BIT_WIDTH_1 = 1;
defparam dpb_inst_7.BLK_SEL_0 = 3'b000;
defparam dpb_inst_7.BLK_SEL_1 = 3'b000;
defparam dpb_inst_7.RESET_MODE = "SYNC";
defparam dpb_inst_7.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFD4BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFC97FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFC87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFC87F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_06 = 256'h0000FFFFFFFFFFFFFDA8FF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_07 = 256'h0000FFFFFFFFFFFC03B17F4FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_08 = 256'h0000FFFFFFFFFFFC00F5FE53FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_09 = 256'h0000FFFFFFFFFFFE0975FE59FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0A = 256'h0000FFFFFFFFFFFE09E5FE007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0B = 256'h0000FFFFFFFFFFFC0AE57E203FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0C = 256'h0000FFFFFFFFFFFC13C2FE401FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0D = 256'h0000FFFFFFFFFFF80BEBFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0E = 256'h0000FFFFFFFFFFF80946FC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0F = 256'h0000FFFFFFFFFFF803C7FC0000FC2940FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_10 = 256'h0000FFFFFFFFFFF817C6FC000079165311940C85FFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_11 = 256'h0000FFFFFFFFFFF023D7FC00007810000000074D52D6CF57FFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_12 = 256'h0000FFFFFFFFFFF00F9FF800007942000000000000000017AAB7FFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_13 = 256'h0000FFFFFFFFFFE00BAFF8100172A0000000000000000000000017FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_14 = 256'h0000FFFFFFFFFFE04BAFF80000F200000000000000000000000017FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_15 = 256'h0000FFFFFFFFFFE08B9FF40001F540000000000000000000000017FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_16 = 256'h0000FFFFFFFFFFC08F8FF00011F520000399C00000000000000016FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_17 = 256'h0000FFFFFFFFFFC08FAFF82000F520000290880300400000000015FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_18 = 256'h0000FFFFFFFFFFC0BE7FE80001F140004310884000A1215000001BFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_19 = 256'h0000FFFFFFFFFF81AF3FE00001F9400207118E8714552A8040000D7FFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_1A = 256'h0000FFFFFFFFFF817FBFE04001E4500140998EC045514A1000000FFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_1B = 256'h0000FFFFFFFFFF811EBFE00003E84000101980605FF94A1481000FBFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_1C = 256'h0000FFFFFFFFFF033EBFC40003EA40004019DE671FF7285FFCA00EFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_1D = 256'h0000FFFFFFFFFF025D5FD40007E5400008119C291FF64508AE200EBFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_1E = 256'h0000FFFFFFFFFE007DBFD40003E1000004304EE21FF6A12806840EBFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_1F = 256'h0000FFFFFFFFFF047DBFFC0447F50000003141064FF6A8DEAE800EBFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_20 = 256'h0000FFFFFFFFFE047BFFFC0E03E10000003184104FFEA2CCAEA00B7FFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_21 = 256'h0000FFFFFFFFFE057BFFAC0407ED8000003108664FF6A22A0E9007FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_22 = 256'h0000FFFFFFFFFE03F3FFA31403DAA00000219C000FF680AA068006BFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_23 = 256'h0000FFFFFFFFFC08F3FF650007F5A00000380C004FF65054560007FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_24 = 256'h0000FFFFFFFFF80975FF290007CA200000318C202FFC7FFFFE0006BFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_25 = 256'h0000FFFFFFFFF809F7FF500017C02000000100E600408001000006BFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_26 = 256'h0000FFFFFFFFF803F7FFD0100FD550000001C06000000000000005DFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_27 = 256'h0000FFFFFFFFF803EBFED0007F93400000000070000402000000077FFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_28 = 256'h0000FFFFFFFFF811EBFE5000FF9510000000000000000090000003FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_29 = 256'h0000FFFFFFFFF007DBFEA580FF95A40000000000000004400000035FFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_2A = 256'h0000FFFFFFFFF007D7FFA2C01FD82A312F80000000000000000003FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_2B = 256'h0000FFFFFFFFF017D7FDE5820FDA0179B42EB72AAABFA800000003FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_2C = 256'h0000FFFFFFFFC01FB7FD58001F5C00000000155717D6AF7F557F7FFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_2D = 256'h0000FFFFFFFF00CFBFFE62021F4A000000000D5E42EFC0000017FBDFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_2E = 256'h0000FFFFFFFF00AFBFFB6A805FD4000000000CD412EF8000000003FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_2F = 256'h0000FFFFFFFF809F5FF9FE801F50000000000D3602E74000000003FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_30 = 256'h0000FFFFFFFFE09F3FFCDE91FF54000000000DB612DA8000000001FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_31 = 256'h0000FFFFFFFFE03FBFBF55D3FF54000000000DFC02FE8000000001B7FFFFFFFF;
defparam dpb_inst_7.INIT_RAM_32 = 256'h0000FFFFFFFFF01F5FFFD393FE58000000000A767FB5C000000001B7FFFFFFFF;
defparam dpb_inst_7.INIT_RAM_33 = 256'h0000FFFFFFFFF82EEFFFE323FE68000000000BD46F754000000001D7FFFFFFFF;
defparam dpb_inst_7.INIT_RAM_34 = 256'h0000FFFFFFFFFC17EFFFFAD3FE68000000000AA46ECB4000000001F7FFFFFFFF;
defparam dpb_inst_7.INIT_RAM_35 = 256'h0000FFFFFFFFFC07F7FFFF27FE68000000000A647FDA4000000001FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_36 = 256'h0000FFFFFFFFFE0BFBFFFF87FE60000000000AF402DFC000000001DFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_37 = 256'h0000FFFFFFFFFE01FBFFFFE7FE68000000000B56ABEEC000000000AFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_38 = 256'h0000FFFFFFFFFF01FDFFFFFFFD6800000000097A0B57C000000000AFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_39 = 256'h0000FFFFFFFFFFC0FEFFFFFFFE70000000001C5C03D6C000000000AFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_3A = 256'h0000FFFFFFFFFFE07FFFFFFFFFF8000000001DD603FE4000000000AFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_3B = 256'h0000FFFFFFFFFFE03F7FFFFFF9D0A51F5152D4E600B54000000000AFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_3C = 256'h0000FFFFFFFFFFF03BBFFFFFFF48F695C4E43D3A355F55F6FA0000EFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_3D = 256'h0000FFFFFFFFFFF81BFFFFFFFFFFFFFFFFFFFFFFFEACA3D6BAD7ABFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_3E = 256'h0000FFFFFFFFFFF80FDFFFFFFFFFFFFFFFFFFFFFFEFFF7FFFDBAEBFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_3F = 256'h0000FFFFFFFFFFFC07EFFFFFFFFFFFFFFFFFFFFFFDDF7AAABEAD5FFFFFFFFFFF;

DPB dpb_inst_8 (
    .DOA({dpb_inst_8_douta_w[14:0],dpb_inst_8_douta[7]}),
    .DOB({dpb_inst_8_doutb_w[14:0],dpb_inst_8_doutb[7]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7]})
);

defparam dpb_inst_8.READ_MODE0 = 1'b1;
defparam dpb_inst_8.READ_MODE1 = 1'b1;
defparam dpb_inst_8.WRITE_MODE0 = 2'b00;
defparam dpb_inst_8.WRITE_MODE1 = 2'b00;
defparam dpb_inst_8.BIT_WIDTH_0 = 1;
defparam dpb_inst_8.BIT_WIDTH_1 = 1;
defparam dpb_inst_8.BLK_SEL_0 = 3'b000;
defparam dpb_inst_8.BLK_SEL_1 = 3'b000;
defparam dpb_inst_8.RESET_MODE = "SYNC";
defparam dpb_inst_8.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFC07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFF07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFF2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFF2FF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_06 = 256'h0000FFFFFFFFFFFFFAF37F1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_07 = 256'h0000FFFFFFFFFFFC046AFE4FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_08 = 256'h0000FFFFFFFFFFFC06A1FEA3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_09 = 256'h0000FFFFFFFFFFFC05D2FEA1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0A = 256'h0000FFFFFFFFFFFE04B3FEA07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0B = 256'h0000FFFFFFFFFFFE01A3FE803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0C = 256'h0000FFFFFFFFFFFC14EBFD001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0D = 256'h0000FFFFFFFFFFFC12E5FC0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0E = 256'h0000FFFFFFFFFFFC13EBFC0003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0F = 256'h0000FFFFFFFFFFF835DAFC0800FD5217FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_10 = 256'h0000FFFFFFFFFFF0235BFE0000FE40A4AA60A05FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_11 = 256'h0000FFFFFFFFFFF816DBFA0000FEC000000010B2AD2830BFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_12 = 256'h0000FFFFFFFFFFF065D7F800007A100000000000000001EAF7DD5FFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_13 = 256'h0000FFFFFFFFFFF06797F810017C0100000000000000000000001BFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_14 = 256'h0000FFFFFFFFFFE057B7F800007D4000000000000000000000001DFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_15 = 256'h0000FFFFFFFFFFE05F6FF00001F00000000000000000000000001DFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_16 = 256'h0000FFFFFFFFFFE02F7FF00011F24000019800000000000000001DFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_17 = 256'h0000FFFFFFFFFFC05B7FF02000FA4000028080470800000000001BFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_18 = 256'h0000FFFFFFFFFFC08FAFE80001ECA0040B38C0675400000000000EFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_19 = 256'h0000FFFFFFFFFFC01EEFE00001E4200087298E664288442800000BFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_1A = 256'h0000FFFFFFFFFF8016DFE04001EA8040023094E0AA04A54548000AFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_1B = 256'h0000FFFFFFFFFF407EBFC80001E200408431A6E92FF2116254000AFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_1C = 256'h0000FFFFFFFFFF805CBFD80007E5000208110C4F4FF783FFFE000BFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_1D = 256'h0000FFFFFFFFFF007D7FD40007D2400200118E654FF690520E000BFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_1E = 256'h0000FFFFFFFFFF015D7FC80007D4C0004011DCEA4FF60A92AE100BFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_1F = 256'h0000FFFFFFFFFE02B97FC40447C0800008188006AFF601CC16200BFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_20 = 256'h0000FFFFFFFFFE02F97F840603CA4000003198800FF6088E06000EFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_21 = 256'h0000FFFFFFFFFE02FA7FA40C07C22000003188470FF60880A6000DDFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_22 = 256'h0000FFFFFFFFFC08FAFFB89C07C5000000138870AFF62400961005FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_23 = 256'h0000FFFFFFFFFC0BFEBF990007C2000000119C050FF6A501068006BFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_24 = 256'h0000FFFFFFFFFC05F6FF540007A18000003184E00FFFFFFFFE8007FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_25 = 256'h0000FFFFFFFFFC13F6FF280017AB800000010047000A1200040007FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_26 = 256'h0000FFFFFFFFF812EDFF200007822000000180E0909020240000077FFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_27 = 256'h0000FFFFFFFFF015EFFE30027FAC1000000000E004000000000007DFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_28 = 256'h0000FFFFFFFFF027EFFEB000FFA1480000000000000004000000055FFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_29 = 256'h0000FFFFFFFFF023EFFEAE00FF6850000000000020000000000007FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_2A = 256'h0000FFFFFFFFF057DBFC4DC01F27D5CEF8000000000000000000037FFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_2B = 256'h0000FFFFFFFFE06BDFFD07820F00D6CE4BF5C8FFFFEA8000000003DFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_2C = 256'h0000FFFFFFFFE047DFFD50001F20000000001EBAFEADDAD5FFD5FDDFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_2D = 256'h0000FFFFFFFF000FAFF9AA021F50000000000AF543BAC00005FFEF7FFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_2E = 256'h0000FFFFFFFF001BAFFA9A801E20000000000BAA13B540000000035FFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_2F = 256'h0000FFFFFFFF800F2FFA1E801F2C000000000BCC03BA8000000002B7FFFFFFFF;
defparam dpb_inst_8.INIT_RAM_30 = 256'h0000FFFFFFFFC0ABFDFD3611FEA4000000000ADC53ADC0000000035FFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_31 = 256'h0000FFFFFFFFE07BBFFF2C43FEA0000010000A5603AB4000000001FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_32 = 256'h0000FFFFFFFFE05FDFFF8C13FEA4000000000B9A7EEA8000000001FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_33 = 256'h0000FFFFFFFFF00FDFFFF403FE90000000000C2E66DFC000000001FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_34 = 256'h0000FFFFFFFFF807EFFFF907FD90000000000D7E67B680000000015FFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_35 = 256'h0000FFFFFFFFFC17F7FFFE53FD90000000000DBE7EB7C00000000157FFFFFFFF;
defparam dpb_inst_8.INIT_RAM_36 = 256'h0000FFFFFFFFFE0BDBFFFF87FD88000000000D9E036AC00000000177FFFFFFFF;
defparam dpb_inst_8.INIT_RAM_37 = 256'h0000FFFFFFFFFF03FBFFFFE7FD90000000000DAA02BB8000000001FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_38 = 256'h0000FFFFFFFFFF81FDFFFFFFFE800000000016D60BFD4000000000FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_39 = 256'h0000FFFFFFFFFF80FEFFFFFFFD800000000017A60B7DC000000000FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_3A = 256'h0000FFFFFFFFFFC0F6FFFFFFFC0400000000122A82ABC000000000FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_3B = 256'h0000FFFFFFFFFFE07B7FFFFFFE2F5AE0AEAFAB5C1DEBC000000000FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_3C = 256'h0000FFFFFFFFFFE83FBFFFFFF4B709EABB5BE2EFDBA9FF5F800000BFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_3D = 256'h0000FFFFFFFFFFF03F9FFFFFFFFFFFFFFFFFFFFAA3535F2D55AADEAFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_3E = 256'h0000FFFFFFFFFFFC0FDFFFFFFFFFFFFFFFFFFFFFBFDBDEEAAFFFDFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_3F = 256'h0000FFFFFFFFFFFE0FEFFFFFFFFFFFFFFFFFFFFFFFFBEFFFD5F7FFFFFFFFFFFF;

DPB dpb_inst_9 (
    .DOA({dpb_inst_9_douta_w[11:0],dpb_inst_9_douta[7:4]}),
    .DOB({dpb_inst_9_doutb_w[11:0],dpb_inst_9_doutb[7:4]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[14],ada[13],ada[12]}),
    .BLKSELB({adb[14],adb[13],adb[12]}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7:4]})
);

defparam dpb_inst_9.READ_MODE0 = 1'b1;
defparam dpb_inst_9.READ_MODE1 = 1'b1;
defparam dpb_inst_9.WRITE_MODE0 = 2'b00;
defparam dpb_inst_9.WRITE_MODE1 = 2'b00;
defparam dpb_inst_9.BIT_WIDTH_0 = 4;
defparam dpb_inst_9.BIT_WIDTH_1 = 4;
defparam dpb_inst_9.BLK_SEL_0 = 3'b100;
defparam dpb_inst_9.BLK_SEL_1 = 3'b100;
defparam dpb_inst_9.RESET_MODE = "SYNC";
defparam dpb_inst_9.INIT_RAM_00 = 256'h7E5F5F5F5F5F5FA7AFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFF7FFEF7FFDFFDFF7FBEFBFD7DFAFE7E;
defparam dpb_inst_9.INIT_RAM_02 = 256'h00000EFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_03 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1;
defparam dpb_inst_9.INIT_RAM_04 = 256'hD7D7D6FA7E5E7EBEFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFF7FEFFBFEFBEFDFBFDF6FAF6FAF6;
defparam dpb_inst_9.INIT_RAM_06 = 256'h100000FFFFFFF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_07 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_08 = 256'h7DF5F6D7D6FAFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFF7FFDFFFDF7FDF7FBEFDFE7E7DFD7DFD;
defparam dpb_inst_9.INIT_RAM_0A = 256'hF00000AFFFFFF2EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_0B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_0C = 256'h7DFDFDFBEBEBEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFEFFEFBFE7FEBFD7EBFBEBEBEBEF;
defparam dpb_inst_9.INIT_RAM_0E = 256'hF5200005FFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_0F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_10 = 256'hF5FD7DF5FDFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFBFF6FF7EF7DF6FDF5FDFDFD7D;
defparam dpb_inst_9.INIT_RAM_12 = 256'hFF500000DFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_13 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_14 = 256'hBFBDF5FAFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFEFFBFFFE7FBFD7EBEBE7DFBFAFBF;
defparam dpb_inst_9.INIT_RAM_16 = 256'hFFF500000FFFFFFF0FFFFFFFFFBFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_17 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_18 = 256'h7F5FBFBFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFDFFFFDF7FBEFBFDFD7DFBFBF6D7FDFD;
defparam dpb_inst_9.INIT_RAM_1A = 256'hFFFF100000EFFFFF7CFFFFFFE7FFFF7FFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1C = 256'hEBE7DFDADBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFEFFFBFFDFFEBFFBFFDFBFBFBFAFBFAF6B;
defparam dpb_inst_9.INIT_RAM_1E = 256'hFFFFF000000FFFFFF1FFFFFFFBFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_20 = 256'h5FBFFA56FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFF7FEFBFE7FBFDFDFBF6FDF6FD7D7DFBFDF;
defparam dpb_inst_9.INIT_RAM_22 = 256'hFFFFFF000000FFFFFF0FFFE7FFBFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_23 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_24 = 256'hBFFE6DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFDF7FD7FFBF7EFAFFBEFD7ED7D7D7D7DE;
defparam dpb_inst_9.INIT_RAM_26 = 256'hFFFFFFF510000CFFFFF0FFE7FEFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_27 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_28 = 256'hFE5DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFDFFBFFBFE7DFBF6F6F5F6F5F6F5F6F5F6F;
defparam dpb_inst_9.INIT_RAM_2A = 256'hFFFFFFFFF10000FFFFD78FFDF7FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2C = 256'hEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFBFEFFBFEBFFBF6FDFBFAF7DF5F5FDBFBFBFBF;
defparam dpb_inst_9.INIT_RAM_2E = 256'hFFFFFFFFFF10000FFFBE5AFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_30 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_31 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFDF7EFDFBFDFDFBF6F5FAF7EBFAFBDF5F5F5F7;
defparam dpb_inst_9.INIT_RAM_32 = 256'hFFFFFFFFFF700000FF5FF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_33 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_35 = 256'hFFFFFFFFFFFFFFFFFFFFFFFDFFBFFBFDFBE7EBF7D7D7DFBEBFAFBDF5F6FAF7FF;
defparam dpb_inst_9.INIT_RAM_36 = 256'hFFFFFFFFFFFF32101EFEBF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_37 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ada[14]),
  .CLK(clka),
  .CE(cea_w)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(dff_q_0),
  .CLK(clka),
  .CE(ocea)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb_w)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(dff_q_2),
  .CLK(clkb),
  .CE(oceb)
);
MUX2 mux_inst_4 (
  .O(douta[0]),
  .I0(dpb_inst_0_douta[0]),
  .I1(dpb_inst_4_douta[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_9 (
  .O(douta[1]),
  .I0(dpb_inst_1_douta[1]),
  .I1(dpb_inst_4_douta[1]),
  .S0(dff_q_1)
);
MUX2 mux_inst_14 (
  .O(douta[2]),
  .I0(dpb_inst_2_douta[2]),
  .I1(dpb_inst_4_douta[2]),
  .S0(dff_q_1)
);
MUX2 mux_inst_19 (
  .O(douta[3]),
  .I0(dpb_inst_3_douta[3]),
  .I1(dpb_inst_4_douta[3]),
  .S0(dff_q_1)
);
MUX2 mux_inst_24 (
  .O(douta[4]),
  .I0(dpb_inst_5_douta[4]),
  .I1(dpb_inst_9_douta[4]),
  .S0(dff_q_1)
);
MUX2 mux_inst_29 (
  .O(douta[5]),
  .I0(dpb_inst_6_douta[5]),
  .I1(dpb_inst_9_douta[5]),
  .S0(dff_q_1)
);
MUX2 mux_inst_34 (
  .O(douta[6]),
  .I0(dpb_inst_7_douta[6]),
  .I1(dpb_inst_9_douta[6]),
  .S0(dff_q_1)
);
MUX2 mux_inst_39 (
  .O(douta[7]),
  .I0(dpb_inst_8_douta[7]),
  .I1(dpb_inst_9_douta[7]),
  .S0(dff_q_1)
);
MUX2 mux_inst_44 (
  .O(doutb[0]),
  .I0(dpb_inst_0_doutb[0]),
  .I1(dpb_inst_4_doutb[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_49 (
  .O(doutb[1]),
  .I0(dpb_inst_1_doutb[1]),
  .I1(dpb_inst_4_doutb[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_54 (
  .O(doutb[2]),
  .I0(dpb_inst_2_doutb[2]),
  .I1(dpb_inst_4_doutb[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_59 (
  .O(doutb[3]),
  .I0(dpb_inst_3_doutb[3]),
  .I1(dpb_inst_4_doutb[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_64 (
  .O(doutb[4]),
  .I0(dpb_inst_5_doutb[4]),
  .I1(dpb_inst_9_doutb[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_69 (
  .O(doutb[5]),
  .I0(dpb_inst_6_doutb[5]),
  .I1(dpb_inst_9_doutb[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_74 (
  .O(doutb[6]),
  .I0(dpb_inst_7_doutb[6]),
  .I1(dpb_inst_9_doutb[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_79 (
  .O(doutb[7]),
  .I0(dpb_inst_8_doutb[7]),
  .I1(dpb_inst_9_doutb[7]),
  .S0(dff_q_3)
);
endmodule //blk_mem_gen_6
