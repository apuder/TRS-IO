//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.05
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9C
//Created Time: Wed Jun 08 05:15:47 2022

module blk_mem_gen_4 (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [5:0] douta;
output [5:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [13:0] ada;
input [5:0] dina;
input [13:0] adb;
input [5:0] dinb;

wire [14:0] dpb_inst_0_douta_w;
wire [14:0] dpb_inst_0_doutb_w;
wire [14:0] dpb_inst_1_douta_w;
wire [14:0] dpb_inst_1_doutb_w;
wire [14:0] dpb_inst_2_douta_w;
wire [14:0] dpb_inst_2_doutb_w;
wire [14:0] dpb_inst_3_douta_w;
wire [14:0] dpb_inst_3_doutb_w;
wire [14:0] dpb_inst_4_douta_w;
wire [14:0] dpb_inst_4_doutb_w;
wire [14:0] dpb_inst_5_douta_w;
wire [14:0] dpb_inst_5_doutb_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[14:0],douta[0]}),
    .DOB({dpb_inst_0_doutb_w[14:0],doutb[0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[0]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b1;
defparam dpb_inst_0.READ_MODE1 = 1'b1;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 1;
defparam dpb_inst_0.BIT_WIDTH_1 = 1;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'hFFFC00000000FFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_01 = 256'hFFD7FFFC00001FFFFFF7FFFC00002FFFFFF7FFF800070FFFFFFFFFFFFC001FFF;
defparam dpb_inst_0.INIT_RAM_02 = 256'hFFE00280000017FFFFE8000000001FFFFFEFFFFE00001FFFFFD79FFE00001FFF;
defparam dpb_inst_0.INIT_RAM_03 = 256'hFFE00000007FCFFFFFE00000FFA00FFFFFEFFFFFC0000FFFFFE9C000000007FF;
defparam dpb_inst_0.INIT_RAM_04 = 256'hFFE0800078000FFFFFE0000000000FFFFFE0000000000FFFFFE0000000000FFF;
defparam dpb_inst_0.INIT_RAM_05 = 256'hFFE000FFFFFE0FFFFFE0007FFFFE0FFFFFE0003FFFF80FFFFFE00007FFE00FFF;
defparam dpb_inst_0.INIT_RAM_06 = 256'hFFE001FFFFFF0FFFFFE001FFFFFF0FFFFFE080FFFFFF0FFFFFE000FFFFFF0FFF;
defparam dpb_inst_0.INIT_RAM_07 = 256'hFFE001FFFFFF0FFFFFE001FFFFFF0FFFFFE001FFFFFF0FFFFFE001FFFFFF0FFF;
defparam dpb_inst_0.INIT_RAM_08 = 256'hFFE001FFFFFF0FFFFFE011FFFFFF0FFFFFE001FFFFFF0FFFFFE001FFFFFF0FFF;
defparam dpb_inst_0.INIT_RAM_09 = 256'hFFE031EFE7FF0FFFFFE3F1FFFFFF0FFFFFE001FFFFFF0FFFFFE001FFFFFF0FFF;
defparam dpb_inst_0.INIT_RAM_0A = 256'hFFE011AAE10307FFFFE011D6EA9B07FFFFE011C6E20307FFFFE011C6E6030FFF;
defparam dpb_inst_0.INIT_RAM_0B = 256'hFFE0119290A707FFFFE01192F0A707FFFFE03192F0A707FFFFE1F182E00307FF;
defparam dpb_inst_0.INIT_RAM_0C = 256'hFFE3F192A62717FFFFE3F19A852717FFFFE0119AC42717FFFFE0119A88A707FF;
defparam dpb_inst_0.INIT_RAM_0D = 256'hFFE031EAE1A717FFFFE3F182E32717FFFFE3F192F22717FFFFE3B192EE2717FF;
defparam dpb_inst_0.INIT_RAM_0E = 256'hFFE011EFF7FF17FFFFE011C6E0A717FFFFE011C6E0A717FFFFE011D6E8A717FF;
defparam dpb_inst_0.INIT_RAM_0F = 256'hFFE0D1FFFFFF17FFFFE011FFFFFF17FFFFE011FFFFFF17FFFFE091FFFFFF17FF;
defparam dpb_inst_0.INIT_RAM_10 = 256'hFFE011FFFFFF17FFFFE011FFFFFF17FFFFE011FFFFFF17FFFFE011FFFFFF17FF;
defparam dpb_inst_0.INIT_RAM_11 = 256'hFFE001FFFFFF17FFFFE001FFFFFF17FFFFE3F1FFFFFF17FFFFE011FFFFFF17FF;
defparam dpb_inst_0.INIT_RAM_12 = 256'hFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FF;
defparam dpb_inst_0.INIT_RAM_13 = 256'hFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FF;
defparam dpb_inst_0.INIT_RAM_14 = 256'hFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FF;
defparam dpb_inst_0.INIT_RAM_15 = 256'hFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FF;
defparam dpb_inst_0.INIT_RAM_16 = 256'hFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FF;
defparam dpb_inst_0.INIT_RAM_17 = 256'hFFE000FFFFFE1FFFFFE000FFFFFE1FFFFFE000FFFFFE1FFFFFE000FFFFFF1FFF;
defparam dpb_inst_0.INIT_RAM_18 = 256'hFFE00003FF811FFFFFE0001FFFE11FFFFFE0003FFFF81FFFFFE0007FFFFC1FFF;
defparam dpb_inst_0.INIT_RAM_19 = 256'hFFE0008000009FFFFFE0000000009FFFFFE0000000001FFFFFE0000000011FFF;
defparam dpb_inst_0.INIT_RAM_1A = 256'hFFE0000000001FFFFFE0000000001FFFFFE0000000001FFFFFE0000B80001FFF;
defparam dpb_inst_0.INIT_RAM_1B = 256'hFFFFFFFFD0003FFFFFF0000000001FFFFFF0000000001FFFFFE0000000001FFF;
defparam dpb_inst_0.INIT_RAM_1C = 256'hFFFFEF85550BFFFFFFFFFF85550BFFFFFFFFFFB555FFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_1D = 256'hFFFF2F81540BFFFFFFFF2F81540BFFFFFFFFAF81540BFFFFFFFF7F81550BFFFF;
defparam dpb_inst_0.INIT_RAM_1E = 256'hFF000000000001FFFFFFFF81540BFFFFFFFFFF81540BFFFFFFFFFF81540BFFFF;
defparam dpb_inst_0.INIT_RAM_1F = 256'hFEFFFFFFFFFFFFFFFEFFFFFFFFFFFEFFFEFFFFFFFFFFFEFFFFFFFFFFFFFFFEFF;
defparam dpb_inst_0.INIT_RAM_20 = 256'hFF800310081403FFFF80003A5C1403FFFF800002FC0003FFFE80001FD00003FF;
defparam dpb_inst_0.INIT_RAM_21 = 256'hFF800000000001FFFF828800000001FFFF838800000001FFFF808010080003FF;
defparam dpb_inst_0.INIT_RAM_22 = 256'hFF1080200020017FFF0000000000017FFF0004281020117FFF801028002011FF;
defparam dpb_inst_0.INIT_RAM_23 = 256'hFD0003E0000001FFFD000FE2050A01FFFF0011C0000001FFFF108000000001FF;
defparam dpb_inst_0.INIT_RAM_24 = 256'hFF0001C10A1011FFFF0003E1000001FFFF0003E0000801FFFD1003E0000801FF;
defparam dpb_inst_0.INIT_RAM_25 = 256'hFF300000000000BFFF300000000000BFFF300000001080FFFF000040000000FF;
defparam dpb_inst_0.INIT_RAM_26 = 256'hFF000000000000FFFF300000000000FFFF300000000000FFFF300000000000BF;
defparam dpb_inst_0.INIT_RAM_27 = 256'hFA2000000FFFFCFFFA007FFC000000FFFE000000000000FFFE000000000000FF;
defparam dpb_inst_0.INIT_RAM_28 = 256'hFFFFFE80000001FFFF000000000000FFFE000000000000FFFA000000000000FF;
defparam dpb_inst_0.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFDF;
defparam dpb_inst_0.INIT_RAM_2A = 256'hF83FFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_2B = 256'hF80083FFFFFFFD1FF8000485F2F1581FF80000000000101FF80000000000001F;
defparam dpb_inst_0.INIT_RAM_2C = 256'hF8000000001FFFDFF80000000000001FF810FFFFFFFFFF5FF8010FFFFFFFFFDF;
defparam dpb_inst_0.INIT_RAM_2D = 256'hF8FFFFFFFFFFFFFFF86FFFFFFFFFFFFFF803FFFFFFFFFFFFF80FFFFFFFFFFFDF;
defparam dpb_inst_0.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000003F;
defparam dpb_inst_0.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DPB dpb_inst_1 (
    .DOA({dpb_inst_1_douta_w[14:0],douta[1]}),
    .DOB({dpb_inst_1_doutb_w[14:0],doutb[1]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[1]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[1]})
);

defparam dpb_inst_1.READ_MODE0 = 1'b1;
defparam dpb_inst_1.READ_MODE1 = 1'b1;
defparam dpb_inst_1.WRITE_MODE0 = 2'b00;
defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
defparam dpb_inst_1.BIT_WIDTH_0 = 1;
defparam dpb_inst_1.BIT_WIDTH_1 = 1;
defparam dpb_inst_1.BLK_SEL_0 = 3'b000;
defparam dpb_inst_1.BLK_SEL_1 = 3'b000;
defparam dpb_inst_1.RESET_MODE = "SYNC";
defparam dpb_inst_1.INIT_RAM_00 = 256'hFFEC00000000FFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_01 = 256'hFFF7FFFC00001FFFFFF7FFFC00001FFFFFF7FFFC00074FFFFFFFFFFFFC000FFF;
defparam dpb_inst_1.INIT_RAM_02 = 256'hFFE00200000007FFFFE80000000017FFFFD7FFFF00001FFFFFD79FFF00001FFF;
defparam dpb_inst_1.INIT_RAM_03 = 256'hFFE00000007FCFFFFFE00000FF800FFFFFE7FFFFC0000FFFFFE1E00000000FFF;
defparam dpb_inst_1.INIT_RAM_04 = 256'hFFE0800078000FFFFFE0000000000FFFFFE0000000000FFFFFE0000000000FFF;
defparam dpb_inst_1.INIT_RAM_05 = 256'hFFE000FFFFFE0FFFFFE0007FFFFE0FFFFFE0003FFFF80FFFFFE00007FFE00FFF;
defparam dpb_inst_1.INIT_RAM_06 = 256'hFFE001FFFFFF0FFFFFE0C0FFFFFF0FFFFFE000FFFFFF0FFFFFE000FFFFFF0FFF;
defparam dpb_inst_1.INIT_RAM_07 = 256'hFFE001FFFFFF0FFFFFE001FFFFFF0FFFFFE001FFFFFF0FFFFFE001FFFFFF0FFF;
defparam dpb_inst_1.INIT_RAM_08 = 256'hFFE001FFFFFF0FFFFFE011FFFFFF0FFFFFE001FFFFFF0FFFFFE001FFFFFF0FFF;
defparam dpb_inst_1.INIT_RAM_09 = 256'hFFE031EFF7FF8FFFFFE3F1FFFFFF8FFFFFE001FFFFFF0FFFFFE001FFFFFF0FFF;
defparam dpb_inst_1.INIT_RAM_0A = 256'hFFE001CBE2638FFFFFE001D3EAFB8FFFFFE001C6E2238FFFFFE001C6E2238FFF;
defparam dpb_inst_1.INIT_RAM_0B = 256'hFFE0019F90E78FFFFFE00193F0E78FFFFFE02193F0E78FFFFFE161A3E3638FFF;
defparam dpb_inst_1.INIT_RAM_0C = 256'hFFE3F19F86678FFFFFE3F19F87678FFFFFE0019FC4678FFFFFE0019F88E78FFF;
defparam dpb_inst_1.INIT_RAM_0D = 256'hFFE031CBE3E78FFFFFE3F1E3E2678FFFFFE3F183E6678FFFFFE2B193E6678FFF;
defparam dpb_inst_1.INIT_RAM_0E = 256'hFFE001EFF7FF8FFFFFE001E6F0A78FFFFFE001C6E0A78FFFFFE001D3EBE78FFF;
defparam dpb_inst_1.INIT_RAM_0F = 256'hFFE041FFFFFF8FFFFFE001FFFFFF8FFFFFE001FFFFFF8FFFFFE0C1FFFFFF8FFF;
defparam dpb_inst_1.INIT_RAM_10 = 256'hFFE001FFFFFF8FFFFFE001FFFFFF8FFFFFE001FFFFFF8FFFFFE001FFFFFF8FFF;
defparam dpb_inst_1.INIT_RAM_11 = 256'hFFE001FFFFFF8FFFFFE001FFFFFF8FFFFFE3F1FFFFFF8FFFFFE001FFFFFF8FFF;
defparam dpb_inst_1.INIT_RAM_12 = 256'hFFE001FFFFFF0FFFFFE001FFFFFF0FFFFFE001FFFFFF0FFFFFE001FFFFFF8FFF;
defparam dpb_inst_1.INIT_RAM_13 = 256'hFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF1FFFFFE001FFFFFF1FFF;
defparam dpb_inst_1.INIT_RAM_14 = 256'hFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FF;
defparam dpb_inst_1.INIT_RAM_15 = 256'hFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FF;
defparam dpb_inst_1.INIT_RAM_16 = 256'hFFE000FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FFFFE001FFFFFF17FF;
defparam dpb_inst_1.INIT_RAM_17 = 256'hFFE000FFFFFE17FFFFE000FFFFFE17FFFFE000FFFFFF17FFFFE000FFFFFF17FF;
defparam dpb_inst_1.INIT_RAM_18 = 256'hFFE00003FF8117FFFFE0001FFFE117FFFFE0003FFFF817FFFFE0007FFFFC17FF;
defparam dpb_inst_1.INIT_RAM_19 = 256'hFFE00080000097FFFFE00100000097FFFFE00000000097FFFFE00000000117FF;
defparam dpb_inst_1.INIT_RAM_1A = 256'hFFE00000000017FFFFE00000000017FFFFE00000000017FFFFE0000F000017FF;
defparam dpb_inst_1.INIT_RAM_1B = 256'hFFFFFFFFF00037FFFFF80000000017FFFFF00000000017FFFFF00000000017FF;
defparam dpb_inst_1.INIT_RAM_1C = 256'hFFFFFFAA8557F7FFFFFFFFAA8557F7FFFFFFFFAAFD5FF7FFFFFFFFFFFFFFF7FF;
defparam dpb_inst_1.INIT_RAM_1D = 256'hFFFF2FAA0153F7FFFFFF27AA0153F7FFFFFF27AA0157F7FFFFFFAFAA8157F7FF;
defparam dpb_inst_1.INIT_RAM_1E = 256'hFF000000000000FFFFFFFFA80153F7FFFFFFFFAA0153F7FFFFFFBFAA0153F7FF;
defparam dpb_inst_1.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_20 = 256'hFF800150205001FFFE800078701001FFFE80004BFC0003FFFEC0007BC00003FF;
defparam dpb_inst_1.INIT_RAM_21 = 256'hFF8000000000017FFF828800000001FFFF83A000000001FFFF828000201001FF;
defparam dpb_inst_1.INIT_RAM_22 = 256'hFF82A000000401FFFF800000000001FFFF8010A01020417FFF8000201020417F;
defparam dpb_inst_1.INIT_RAM_23 = 256'hFF0001E0000001FFFF0005E0040811FFFF0001E0000001FFFF008020000001FF;
defparam dpb_inst_1.INIT_RAM_24 = 256'hFF0002C4081030FFFD000344000000FFFD1003E0000001FFFD1001E0000201FF;
defparam dpb_inst_1.INIT_RAM_25 = 256'hFF380000000000FFFF180000000000BFFF100000000400BFFF000000000000BF;
defparam dpb_inst_1.INIT_RAM_26 = 256'hFF000000000000FFFF300000000000FFFF300000000000FFFF380000000000FF;
defparam dpb_inst_1.INIT_RAM_27 = 256'hFE3000003FFFFCFFFF007FFA000000FFFF000000000000FFFF000000000000FF;
defparam dpb_inst_1.INIT_RAM_28 = 256'hFBFFFF00000009DFFB000000000000DFFB000000000000FFFE000000000000FF;
defparam dpb_inst_1.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_2A = 256'hF82FFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_2B = 256'hF80087BDFFFFFF3FF800001DF861F81FF80000000000001FF80000000000001F;
defparam dpb_inst_1.INIT_RAM_2C = 256'hF8000000001FFFDFF80000000000001FF805FFFFFFFFFFDFF8000FFFFFFFFFDF;
defparam dpb_inst_1.INIT_RAM_2D = 256'hF8FFFFFFFFFFFFDFF83FFFFFFFFFFFDFF80BFFFFFFFFFFDFF80DFFFFFFFFFFDF;
defparam dpb_inst_1.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000001F;
defparam dpb_inst_1.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DPB dpb_inst_2 (
    .DOA({dpb_inst_2_douta_w[14:0],douta[2]}),
    .DOB({dpb_inst_2_doutb_w[14:0],doutb[2]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[2]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[2]})
);

defparam dpb_inst_2.READ_MODE0 = 1'b1;
defparam dpb_inst_2.READ_MODE1 = 1'b1;
defparam dpb_inst_2.WRITE_MODE0 = 2'b00;
defparam dpb_inst_2.WRITE_MODE1 = 2'b00;
defparam dpb_inst_2.BIT_WIDTH_0 = 1;
defparam dpb_inst_2.BIT_WIDTH_1 = 1;
defparam dpb_inst_2.BLK_SEL_0 = 3'b000;
defparam dpb_inst_2.BLK_SEL_1 = 3'b000;
defparam dpb_inst_2.RESET_MODE = "SYNC";
defparam dpb_inst_2.INIT_RAM_00 = 256'hFFEC00000000FFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_01 = 256'hFFF7FFFE00001FFFFFF7FFFC00001FFFFFFFFFFC00079FFFFFEFFFFFFC000FFF;
defparam dpb_inst_2.INIT_RAM_02 = 256'hFFE0028000000FFFFFD00000000007FFFFD7FFFF000017FFFFF78FFF00001FFF;
defparam dpb_inst_2.INIT_RAM_03 = 256'hFFE00000007FEFFFFFE000007F800FFFFFE7FFFFE0000FFFFFE5800000000FFF;
defparam dpb_inst_2.INIT_RAM_04 = 256'hFFE0000078000FFFFFE0000000000FFFFFE0000000000FFFFFE0000000000FFF;
defparam dpb_inst_2.INIT_RAM_05 = 256'hFFE000FFFFFF0FFFFFE0007FFFFE0FFFFFE0003FFFFC0FFFFFE00007FFE00FFF;
defparam dpb_inst_2.INIT_RAM_06 = 256'hFFE000FFFFFF0FFFFFE040FFFFFF0FFFFFE000FFFFFF0FFFFFE000FFFFFF0FFF;
defparam dpb_inst_2.INIT_RAM_07 = 256'hFFE001FFFFFF8FFFFFE001FFFFFF0FFFFFE001FFFFFF0FFFFFE001FFFFFF0FFF;
defparam dpb_inst_2.INIT_RAM_08 = 256'hFFE001FFFFFF8FFFFFE011FFFFFF8FFFFFE001FFFFFF8FFFFFE001FFFFFF8FFF;
defparam dpb_inst_2.INIT_RAM_09 = 256'hFFE231EFF7FF8FFFFFE3F1FFFFFF8FFFFFE001FFFFFF8FFFFFE001FFFFFF8FFF;
defparam dpb_inst_2.INIT_RAM_0A = 256'hFFE001C2F2638FFFFFE001DAFAFB8FFFFFE001C6F2238FFFFFE001E6F3238FFF;
defparam dpb_inst_2.INIT_RAM_0B = 256'hFFE0019E92F78FFFFFE0019EF3F78FFFFFE0A1E2F3F78FFFFFE1E1E2F3638FFF;
defparam dpb_inst_2.INIT_RAM_0C = 256'hFFE3F19E86F78FFFFFE3F19A86778FFFFFE0019ACB778FFFFFE0019A93F78FFF;
defparam dpb_inst_2.INIT_RAM_0D = 256'hFFE211C2E2778FFFFFE3F1E2E2778FFFFFE3F1E2E6778FFFFFE3319EE6778FFF;
defparam dpb_inst_2.INIT_RAM_0E = 256'hFFE001FFFFFF8FFFFFE001E6F0B78FFFFFE001C6E2B78FFFFFE001D2EF378FFF;
defparam dpb_inst_2.INIT_RAM_0F = 256'hFFE0C1FFFFFF8FFFFFE001FFFFFF8FFFFFE001FFFFFF8FFFFFE0C1FFFFFF8FFF;
defparam dpb_inst_2.INIT_RAM_10 = 256'hFFE001FFFFFF8FFFFFE001FFFFFF8FFFFFE001FFFFFF8FFFFFE001FFFFFF8FFF;
defparam dpb_inst_2.INIT_RAM_11 = 256'hFFE001FFFFFF8FFFFFE001FFFFFF8FFFFFE3F1FFFFFF8FFFFFE201FFFFFF8FFF;
defparam dpb_inst_2.INIT_RAM_12 = 256'hFFE001FFFFFF8FFFFFE001FFFFFF8FFFFFE001FFFFFF8FFFFFE001FFFFFF8FFF;
defparam dpb_inst_2.INIT_RAM_13 = 256'hFFE001FFFFFF8FFFFFE001FFFFFF8FFFFFE001FFFFFF8FFFFFE001FFFFFF8FFF;
defparam dpb_inst_2.INIT_RAM_14 = 256'hFFE001FFFFFF0FFFFFE001FFFFFF0FFFFFE001FFFFFF0FFFFFE001FFFFFF8FFF;
defparam dpb_inst_2.INIT_RAM_15 = 256'hFFE001FFFFFF0FFFFFE001FFFFFF0FFFFFE001FFFFFF0FFFFFE001FFFFFF0FFF;
defparam dpb_inst_2.INIT_RAM_16 = 256'hFFE000FFFFFF0FFFFFE000FFFFFF0FFFFFE000FFFFFF0FFFFFE000FFFFFF0FFF;
defparam dpb_inst_2.INIT_RAM_17 = 256'hFFE000FFFFFE0FFFFFE000FFFFFE0FFFFFE000FFFFFF0FFFFFE000FFFFFF0FFF;
defparam dpb_inst_2.INIT_RAM_18 = 256'hFFE00003FF811FFFFFE0001FFFE11FFFFFE0003FFFFD0FFFFFE0007FFFFE0FFF;
defparam dpb_inst_2.INIT_RAM_19 = 256'hFFE0008000001FFFFFE0000000009FFFFFE0000000009FFFFFE0000000001FFF;
defparam dpb_inst_2.INIT_RAM_1A = 256'hFFF0000000001FFFFFE0000000001FFFFFE0000000001FFFFFE0000B80001FFF;
defparam dpb_inst_2.INIT_RAM_1B = 256'hFFFFFFFFF0003FFFFFF8000000001FFFFFF0000000001FFFFFF0000000001FFF;
defparam dpb_inst_2.INIT_RAM_1C = 256'hFFFFFF82AA07FFFFFFFFFFC2AA87FFFFFFFFFFDAAAFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1D = 256'hFFFFA782AA07F7FFFFFFA782AA07F7FFFFFFE782AA07F7FFFFFFA782AA07F7FF;
defparam dpb_inst_2.INIT_RAM_1E = 256'hFF000000000000FFFFFFFF80A807FFFFFFFFFF80AA07F7FFFFFFAF80AA07F7FF;
defparam dpb_inst_2.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_20 = 256'hFE800140A04021FFFF800061705021FFFF800041FE0001FFFFC0007DC20003FF;
defparam dpb_inst_2.INIT_RAM_21 = 256'hFF801000000001FFFF8204000000017FFE8E00000000017FFE8200002040017F;
defparam dpb_inst_2.INIT_RAM_22 = 256'hFF82A000000001FFFF800000000001FFFF8008A0408141FFFF801020408141FF;
defparam dpb_inst_2.INIT_RAM_23 = 256'hFF0001E0000000FFFF8005E0042811FFFF8001E0000001FFFF828000000009FF;
defparam dpb_inst_2.INIT_RAM_24 = 256'hFD000184281080BFFF000160000000BFFF0081E0000000FFFF0081E0002000FF;
defparam dpb_inst_2.INIT_RAM_25 = 256'hFF180000000000FFFF188000000000FFFD188000000080FFFD000000000000BF;
defparam dpb_inst_2.INIT_RAM_26 = 256'hFF000000000000FFFF180000000000FFFF180000000000FFFF180000000000FF;
defparam dpb_inst_2.INIT_RAM_27 = 256'hFF3800000FFFFE5FFF007FEC0000007FFF000000000000FFFF000000000000FF;
defparam dpb_inst_2.INIT_RAM_28 = 256'hFBFFFF00000004FFFF000000000000FFFF0000000000005FFF0000000000005F;
defparam dpb_inst_2.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFBFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2A = 256'hF80FFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2B = 256'hF80085EFFFFFFC1FF8000083FA74F81FF80000000000001FF80000000000001F;
defparam dpb_inst_2.INIT_RAM_2C = 256'hFC000000000FFFDFFC0000000000001FF807BFFFFFFFFFFFF80027FFFFFFFF9F;
defparam dpb_inst_2.INIT_RAM_2D = 256'hFCFFFFFFFFFFFFDFFC17FFFFFFFFFFFFFC0BFFFFFFFFFFFFFC05FFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000001F;
defparam dpb_inst_2.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DPB dpb_inst_3 (
    .DOA({dpb_inst_3_douta_w[14:0],douta[3]}),
    .DOB({dpb_inst_3_doutb_w[14:0],doutb[3]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[3]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[3]})
);

defparam dpb_inst_3.READ_MODE0 = 1'b1;
defparam dpb_inst_3.READ_MODE1 = 1'b1;
defparam dpb_inst_3.WRITE_MODE0 = 2'b00;
defparam dpb_inst_3.WRITE_MODE1 = 2'b00;
defparam dpb_inst_3.BIT_WIDTH_0 = 1;
defparam dpb_inst_3.BIT_WIDTH_1 = 1;
defparam dpb_inst_3.BLK_SEL_0 = 3'b000;
defparam dpb_inst_3.BLK_SEL_1 = 3'b000;
defparam dpb_inst_3.RESET_MODE = "SYNC";
defparam dpb_inst_3.INIT_RAM_00 = 256'hFFFE000000007FFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_01 = 256'hFFF7FFFE00001FFFFFF3FFFE00001FFFFFEBFFFC0003CFFFFFEFFFFFFE000FFF;
defparam dpb_inst_3.INIT_RAM_02 = 256'hFFF001C000000FFFFFD0000000000FFFFFF7FFFF000017FFFFF79FFF000017FF;
defparam dpb_inst_3.INIT_RAM_03 = 256'hFFF0000000BFEFFFFFF000007FA00FFFFFF7FFFFE0000FFFFFF5C00000000FFF;
defparam dpb_inst_3.INIT_RAM_04 = 256'hFFE0400078000FFFFFE0000000000FFFFFE0000000000FFFFFE0000000000FFF;
defparam dpb_inst_3.INIT_RAM_05 = 256'hFFE0007FFFFF0FFFFFE0007FFFFE0FFFFFE0003FFFFC0FFFFFE00007FFF00FFF;
defparam dpb_inst_3.INIT_RAM_06 = 256'hFFE000FFFFFF0FFFFFE000FFFFFF0FFFFFE040FFFFFF0FFFFFE000FFFFFF0FFF;
defparam dpb_inst_3.INIT_RAM_07 = 256'hFFE000FFFFFF8FFFFFE000FFFFFF8FFFFFE000FFFFFF8FFFFFE000FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_08 = 256'hFFE001FFFFFF8FFFFFE011FFFFFF8FFFFFE001FFFFFF8FFFFFE001FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_09 = 256'hFFE231E7F7FF8FFFFFE3F1FFFFFF8FFFFFE001FFFFFF8FFFFFE001FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_0A = 256'hFFE201C2760B8FFFFFE201DA7ADF8FFFFFE201C272038FFFFFE201E673038FFF;
defparam dpb_inst_3.INIT_RAM_0B = 256'hFFE201D8139F8FFFFFE201FA779F8FFFFFE241E67E9F8FFFFFE3E1C2760B8FFF;
defparam dpb_inst_3.INIT_RAM_0C = 256'hFFE3F1D8069F8FFFFFE3F1D80E1F8FFFFFE20198321F8FFFFFE201D8139F8FFF;
defparam dpb_inst_3.INIT_RAM_0D = 256'hFFE211C2621F8FFFFFC3F1C2621F8FFFFFE3F1E6661F8FFFFFE311FA661F8FFF;
defparam dpb_inst_3.INIT_RAM_0E = 256'hFFC201FFFFFF8FFFFFC201E672978FFFFFE201E272178FFFFFC201DA661F8FFF;
defparam dpb_inst_3.INIT_RAM_0F = 256'hFFE261FFFFFF8FFFFFC281FFFFFF8FFFFFE201FFFFFF8FFFFFC241FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_10 = 256'hFFE201FFFFFF8FFFFFC201FFFFFF8FFFFFC201FFFFFF8FFFFFC201FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_11 = 256'hFFC001FFFFFF8FFFFFC001FFFFFF8FFFFFC3F1FFFFFF8FFFFFC201FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_12 = 256'hFFD001FFFFFF8FFFFFC001FFFFFF8FFFFFC001FFFFFF8FFFFFC001FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_13 = 256'hFFD001FFFFFF8FFFFFD001FFFFFF8FFFFFD001FFFFFF8FFFFFD001FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_14 = 256'hFFD001FFFFFF8FFFFFD001FFFFFF8FFFFFD001FFFFFF8FFFFFD001FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_15 = 256'hFFD000FFFFFF0FFFFFD000FFFFFF0FFFFFD000FFFFFF8FFFFFD001FFFFFF8FFF;
defparam dpb_inst_3.INIT_RAM_16 = 256'hFFD000FFFFFF0FFFFFD000FFFFFF0FFFFFD000FFFFFF0FFFFFD000FFFFFF0FFF;
defparam dpb_inst_3.INIT_RAM_17 = 256'hFFD0007FFFFE0FFFFFD000FFFFFF0FFFFFD000FFFFFF0FFFFFD000FFFFFF0FFF;
defparam dpb_inst_3.INIT_RAM_18 = 256'hFFD00003FF810FFFFFD0000FFFF10FFFFFD0003FFFFC0FFFFFD0007FFFFE0FFF;
defparam dpb_inst_3.INIT_RAM_19 = 256'hFFD0008000000FFFFFD0000000000FFFFFD0000000008FFFFFD0000000008FFF;
defparam dpb_inst_3.INIT_RAM_1A = 256'hFFD0000000000FFFFFD0000000000FFFFFD0000000000FFFFFD0000F80000FFF;
defparam dpb_inst_3.INIT_RAM_1B = 256'hFFDFFFFFF0003FFFFFD8000000001FFFFFD0000000001FFFFFD0000000001FFF;
defparam dpb_inst_3.INIT_RAM_1C = 256'hFFDFFFD502ABFFFFFFDFFFD502ABFFFFFFDFFFD57EBFFFFFFFDFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_1D = 256'hFFDFA7D502ABFFFFFFDFA7D502ABFFFFFFDFAFD502ABFFFFFFDFF7D502ABFFFF;
defparam dpb_inst_3.INIT_RAM_1E = 256'hFF000000000000FFFFDFFFD400A3FFFFFFDFFFD402ABFFFFFFDFF7D402ABFFFF;
defparam dpb_inst_3.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_20 = 256'hFF8001408140817FFF800041C140817FFF800001D60001FFFFC0003FE20003FF;
defparam dpb_inst_3.INIT_RAM_21 = 256'hFE800000000001FFFE8A0000000001FFFE8E0400000001FFFF8800008100817F;
defparam dpb_inst_3.INIT_RAM_22 = 256'hFF8A0030003001FFFF801000003001FFFF801281000101FFFE800001008101FF;
defparam dpb_inst_3.INIT_RAM_23 = 256'hFF8001E0000000FFFF8005E8002040FFFF8001E8000000FFFF820000000001FF;
defparam dpb_inst_3.INIT_RAM_24 = 256'hFF000080204090FFFF0001E0000000FFFF8201E0000400BFFF8201E0000400BF;
defparam dpb_inst_3.INIT_RAM_25 = 256'hFD180000000000FFFD188000000000FFFF188000001800FFFF000000000800FF;
defparam dpb_inst_3.INIT_RAM_26 = 256'hFF0000000000007FFF180000000000FFFF180000000000FFFD180000000000FF;
defparam dpb_inst_3.INIT_RAM_27 = 256'hFF30000037FFFE5FFF007FF80000005FFF0000000000005FFF0000000000007F;
defparam dpb_inst_3.INIT_RAM_28 = 256'hFFFFFE00000004FFFF000000000000FFFF0000000000007FFF0000000000007F;
defparam dpb_inst_3.INIT_RAM_29 = 256'hFBFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2A = 256'hF82FFFFFFFFFFF9FFBFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFBFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2B = 256'hF8000DDFFFFDFC9FF8000081F75DF01FF80000000000001FF80000000000001F;
defparam dpb_inst_3.INIT_RAM_2C = 256'hFC000000001FFFDFFC0000000000001FFC18FFFFFFFFFFFFF8008F3FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2D = 256'hFC7FFFFFFFFFFFFFFC1FFFFFFFFFFFFFFC31FFFFFFFFFFFFFC27FFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000001F;
defparam dpb_inst_3.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DPB dpb_inst_4 (
    .DOA({dpb_inst_4_douta_w[14:0],douta[4]}),
    .DOB({dpb_inst_4_doutb_w[14:0],doutb[4]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[4]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[4]})
);

defparam dpb_inst_4.READ_MODE0 = 1'b1;
defparam dpb_inst_4.READ_MODE1 = 1'b1;
defparam dpb_inst_4.WRITE_MODE0 = 2'b00;
defparam dpb_inst_4.WRITE_MODE1 = 2'b00;
defparam dpb_inst_4.BIT_WIDTH_0 = 1;
defparam dpb_inst_4.BIT_WIDTH_1 = 1;
defparam dpb_inst_4.BLK_SEL_0 = 3'b000;
defparam dpb_inst_4.BLK_SEL_1 = 3'b000;
defparam dpb_inst_4.RESET_MODE = "SYNC";
defparam dpb_inst_4.INIT_RAM_00 = 256'hFFFE000000007FFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_01 = 256'hFFF7FFFE000017FFFFEBFFFE00001FFFFFEBFFFC00038FFFFFFFFFFFFE000FFF;
defparam dpb_inst_4.INIT_RAM_02 = 256'hFFD0018000000FFFFFF0000000000FFFFFF7FFFF00000FFFFFF79FFF000017FF;
defparam dpb_inst_4.INIT_RAM_03 = 256'hFFD00000007FEFFFFFD000003FA00FFFFFD7FFFFE0000BFFFFD1A00000000FFF;
defparam dpb_inst_4.INIT_RAM_04 = 256'hFFD0400078000FFFFFD0000000000FFFFFD0000000000FFFFFD0000000000FFF;
defparam dpb_inst_4.INIT_RAM_05 = 256'hFFD0007FFFFF0FFFFFD0007FFFFE0FFFFFD0003FFFFC0FFFFFD00007FFF00FFF;
defparam dpb_inst_4.INIT_RAM_06 = 256'hFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD040FFFFFF0FFFFFD000FFFFFF0FFF;
defparam dpb_inst_4.INIT_RAM_07 = 256'hFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_08 = 256'hFFD000FFFFFF8FFFFFD010FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_09 = 256'hFFD210F7F7FF8FFFFFD3F0FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_0A = 256'hFFD201C276038FFFFFD201DA76CF8FFFFFD201E273038FFFFFD201E673038FFF;
defparam dpb_inst_4.INIT_RAM_0B = 256'hFFD201F812938FFFFFD201F87E938FFFFFD211C878138FFFFFD3B1C670038FFF;
defparam dpb_inst_4.INIT_RAM_0C = 256'hFFD3F1F81E938FFFFFD3F1F81A138FFFFFD201F832138FFFFFD201F812138FFF;
defparam dpb_inst_4.INIT_RAM_0D = 256'hFFD211D278138FFFFFD3F1C660138FFFFFD3F1C066138FFFFFD331E866938FFF;
defparam dpb_inst_4.INIT_RAM_0E = 256'hFFD201FFFBFF8FFFFFD201E670138FFFFFD201E270138FFFFFD201CA74138FFF;
defparam dpb_inst_4.INIT_RAM_0F = 256'hFFD201FFFFFF8FFFFFD201FFFFFF8FFFFFD201FFFFFF8FFFFFD281FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_10 = 256'hFFD201FFFFFF8FFFFFD201FFFFFF8FFFFFD201FFFFFF8FFFFFD201FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_11 = 256'hFFD001FFFFFF8FFFFFD001FFFFFF8FFFFFD3F1FFFFFF8FFFFFD201FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_12 = 256'hFFD001FFFFFF8FFFFFD001FFFFFF8FFFFFD001FFFFFF8FFFFFD001FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_13 = 256'hFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD001FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_14 = 256'hFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_15 = 256'hFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_16 = 256'hFFD000FFFFFF0FFFFFD000FFFFFF0FFFFFD000FFFFFF8FFFFFD000FFFFFF8FFF;
defparam dpb_inst_4.INIT_RAM_17 = 256'hFFD0007FFFFE0FFFFFD0007FFFFF0FFFFFD000FFFFFF0FFFFFD000FFFFFF0FFF;
defparam dpb_inst_4.INIT_RAM_18 = 256'hFFD00003FF808FFFFFD0000FFFF10FFFFFD0003FFFFC0FFFFFD0007FFFFE0FFF;
defparam dpb_inst_4.INIT_RAM_19 = 256'hFFD0008000000FFFFFD0000000000FFFFFD0000000008FFFFFD0000000008FFF;
defparam dpb_inst_4.INIT_RAM_1A = 256'hFFD0000000000FFFFFD0000000000FFFFFD0000002000FFFFFD0000F80004FFF;
defparam dpb_inst_4.INIT_RAM_1B = 256'hFFDFFFFFF0001FFFFFD8000000001FFFFFD0000000001FFFFFD0000000000FFF;
defparam dpb_inst_4.INIT_RAM_1C = 256'hFFDFF7C1550BFFFFFFDFFFC1550BFFFFFFDFFFED55FFFFFFFFDFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1D = 256'hFFDFB7C1540BFFFFFFDFB7C1550BFFFFFFDFB7C1550BFFFFFFDFF7C1550BFFFF;
defparam dpb_inst_4.INIT_RAM_1E = 256'hFF000000000000FFFFDFFFC0540BFFFFFFDFFFC0540BFFFFFFDFF7C1540BFFFF;
defparam dpb_inst_4.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_20 = 256'hFF800102010081FFFFC000054300817FFFC00001FE00017FFFC0003FE000017F;
defparam dpb_inst_4.INIT_RAM_21 = 256'hFF800000000001FFFF8A0000000001FFFF880000000001FFFF880002010001FF;
defparam dpb_inst_4.INIT_RAM_22 = 256'hFF8A0020001000FFFE800810000000FFFE800A81020501FFFE800001020501FF;
defparam dpb_inst_4.INIT_RAM_23 = 256'hFF8001E0000800BFFF8005E0508140BFFF8001E0000000BFFF8A0000000020FF;
defparam dpb_inst_4.INIT_RAM_24 = 256'hFF8000B0214210FFFF8001F0000000FFFF8201E0000008FFFF8201E0000508FF;
defparam dpb_inst_4.INIT_RAM_25 = 256'hFF180000000000FFFF188000000000FFFF188000000200FFFF800000000800FF;
defparam dpb_inst_4.INIT_RAM_26 = 256'hFD0000000000005FFD1800000000007FFD1800000000007FFD180000000000FF;
defparam dpb_inst_4.INIT_RAM_27 = 256'hFF30000007FFFE7FFF007FF20000007FFF0000000000007FFF0000000000005F;
defparam dpb_inst_4.INIT_RAM_28 = 256'hFFFFFE80000000FFFF0000000000007FFF0000000000007FFF0000000000007F;
defparam dpb_inst_4.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2A = 256'hFC17FFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2B = 256'hFC00065FFFFFFC9FFC000221FF74F81FFC0000000000001FFC0000000000001F;
defparam dpb_inst_4.INIT_RAM_2C = 256'hFC000000001FFFFFFC0000000000001FFC0EFF7FFFFFFFBFFC02876FFFFFFEBF;
defparam dpb_inst_4.INIT_RAM_2D = 256'hFCFFFFFFFFFFFFFFFC6FFFFFFFFFFFFFFC0BFFFFFFFFFFFFFC0FFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000001F;
defparam dpb_inst_4.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DPB dpb_inst_5 (
    .DOA({dpb_inst_5_douta_w[14:0],douta[5]}),
    .DOB({dpb_inst_5_doutb_w[14:0],doutb[5]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,gw_gnd}),
    .BLKSELB({gw_gnd,gw_gnd,gw_gnd}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[5]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[5]})
);

defparam dpb_inst_5.READ_MODE0 = 1'b1;
defparam dpb_inst_5.READ_MODE1 = 1'b1;
defparam dpb_inst_5.WRITE_MODE0 = 2'b00;
defparam dpb_inst_5.WRITE_MODE1 = 2'b00;
defparam dpb_inst_5.BIT_WIDTH_0 = 1;
defparam dpb_inst_5.BIT_WIDTH_1 = 1;
defparam dpb_inst_5.BLK_SEL_0 = 3'b000;
defparam dpb_inst_5.BLK_SEL_1 = 3'b000;
defparam dpb_inst_5.RESET_MODE = "SYNC";
defparam dpb_inst_5.INIT_RAM_00 = 256'hFFFE000000007FFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_01 = 256'hFFEBFFFE000017FFFFEBFFFE000017FFFFFBFFFC00038FFFFFFFFFFFFE000FFF;
defparam dpb_inst_5.INIT_RAM_02 = 256'hFFF001C000000FFFFFF0000000000FFFFFF7EFFF00000FFFFFF7CFFF00000FFF;
defparam dpb_inst_5.INIT_RAM_03 = 256'hFFF00000007FEBFFFFF000007F800BFFFFF7FFFFE0000BFFFFF4C00000000BFF;
defparam dpb_inst_5.INIT_RAM_04 = 256'hFFF040007C000BFFFFF0000000000BFFFFF0000000001BFFFFF0000000000BFF;
defparam dpb_inst_5.INIT_RAM_05 = 256'hFFF0007FFFFF0BFFFFF0003FFFFE0BFFFFF0001FFFFC0BFFFFF00003FFF00BFF;
defparam dpb_inst_5.INIT_RAM_06 = 256'hFFF000FFFFFF8BFFFFF000FFFFFF8BFFFFF040FFFFFF8BFFFFF0007FFFFF0BFF;
defparam dpb_inst_5.INIT_RAM_07 = 256'hFFF000FFFFFF8BFFFFF000FFFFFF8BFFFFF000FFFFFF8BFFFFF000FFFFFF8BFF;
defparam dpb_inst_5.INIT_RAM_08 = 256'hFFF000FFFFFF8BFFFFF010FFFFFF8BFFFFF000FFFFFF8BFFFFF000FFFFFF8BFF;
defparam dpb_inst_5.INIT_RAM_09 = 256'hFFF018F7F3FF8BFFFFF1F0FFFFFF8BFFFFF000FFFFFF8BFFFFF000FFFFFF8BFF;
defparam dpb_inst_5.INIT_RAM_0A = 256'hFFF008D670818BFFFFF008CA744D8BFFFFF008E273018BFFFFF008E273018BFF;
defparam dpb_inst_5.INIT_RAM_0B = 256'hFFF008D814138BFFFFF008C878138BFFFFF038C878138BFFFFF1B8C070018BFF;
defparam dpb_inst_5.INIT_RAM_0C = 256'hFFF1F8D81A938BFFFFF1F8D812138BFFFFF008F832138BFFFFF008D812138BFF;
defparam dpb_inst_5.INIT_RAM_0D = 256'hFFF018D270138FFFFFF1F8C478138FFFFFF1F9C87D938FFFFFF159C87F138BFF;
defparam dpb_inst_5.INIT_RAM_0E = 256'hFFF009F7FBFF8FFFFFF009E270138FFFFFF008E270138FFFFFF008EA74138FFF;
defparam dpb_inst_5.INIT_RAM_0F = 256'hFFF028FFFFFF8FFFFFF009FFFFFF8FFFFFF009FFFFFF8FFFFFF069FFFFFF8FFF;
defparam dpb_inst_5.INIT_RAM_10 = 256'hFFF008FFFFFF8FFFFFF008FFFFFF8FFFFFF008FFFFFF8FFFFFF008FFFFFF8FFF;
defparam dpb_inst_5.INIT_RAM_11 = 256'hFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF1F8FFFFFF8FFFFFF008FFFFFF8FFF;
defparam dpb_inst_5.INIT_RAM_12 = 256'hFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFF;
defparam dpb_inst_5.INIT_RAM_13 = 256'hFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFF;
defparam dpb_inst_5.INIT_RAM_14 = 256'hFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFF;
defparam dpb_inst_5.INIT_RAM_15 = 256'hFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFF;
defparam dpb_inst_5.INIT_RAM_16 = 256'hFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFFFFF000FFFFFF8FFF;
defparam dpb_inst_5.INIT_RAM_17 = 256'hFFF0007FFFFF0FFFFFF0007FFFFF0FFFFFF0007FFFFF0FFFFFF000FFFFFF0FFF;
defparam dpb_inst_5.INIT_RAM_18 = 256'hFFF00001FF808FFFFFF0000FFFF00FFFFFF0001FFFFC0FFFFFF0007FFFFE0FFF;
defparam dpb_inst_5.INIT_RAM_19 = 256'hFFF0008000004FFFFFF0000000000FFFFFF0000000008FFFFFF0000000008FFF;
defparam dpb_inst_5.INIT_RAM_1A = 256'hFFF0000000000FFFFFF0000000000FFFFFF0000000000FFFFFF0000580004FFF;
defparam dpb_inst_5.INIT_RAM_1B = 256'hFFFFFFFFF0001FFFFFF8000000001FFFFFF8000000000FFFFFF0000000000FFF;
defparam dpb_inst_5.INIT_RAM_1C = 256'hFFFFF7EA8157FFFFFFFFFFEA8157FFFFFFFFFFEABD5FFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_1D = 256'hFFFFB7EA0155FFFFFFFFB7EA0155FFFFFFFFB7EA8155FFFFFFFFBFEA8155FFFF;
defparam dpb_inst_5.INIT_RAM_1E = 256'hFF800000000000FFFFFFFFEA0151FFFFFFFFFFEA0151FFFFFFFFFFEA0151FFFF;
defparam dpb_inst_5.INIT_RAM_1F = 256'hFFFFFFFFFFFFFF7FFFFFFFFFFFFFFF7FFF7FFFFFFFFFFFFFFF7FFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_20 = 256'hFFC00102050201FFFFC0000D0F0201FFFFC00005FE0001FFFFC0003FEA00017F;
defparam dpb_inst_5.INIT_RAM_21 = 256'hFF800000000000FFFF880000000001FFFFC84400000001FFFFC04002000201FF;
defparam dpb_inst_5.INIT_RAM_22 = 256'hFE880000000400BFFF800800000000FFFF800A05080400FFFF8010040A0400FF;
defparam dpb_inst_5.INIT_RAM_23 = 256'hFF8001F0000000FFFF800DE0408100FFFE8009E0000000BFFE880000000008BF;
defparam dpb_inst_5.INIT_RAM_24 = 256'hFF8000A0210208FFFF8001B0000000FFFF8201F0000000FFFF8A01F0000000FF;
defparam dpb_inst_5.INIT_RAM_25 = 256'hFF9808000000007FFF980000000000FFFF988000000240FFFF800020000000FF;
defparam dpb_inst_5.INIT_RAM_26 = 256'hFD0000000000007FFF1800000000005FFF1800000000005FFF9800000000007F;
defparam dpb_inst_5.INIT_RAM_27 = 256'hFF30000007FFFE7FFF003FFF0000007FFD0000000000007FFD0000000000007F;
defparam dpb_inst_5.INIT_RAM_28 = 256'hFFFFFF80000006FFFF8000000000007FFF0000000000007FFF0000000000007F;
defparam dpb_inst_5.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_2A = 256'hFC17FFFFFFFFFF0FFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFEF;
defparam dpb_inst_5.INIT_RAM_2B = 256'hFC0003F7FFF7FE9FFC000262FF7DD41FFC0000000000000FFC0000000000000F;
defparam dpb_inst_5.INIT_RAM_2C = 256'hFC000000000FFFFFFC0000000000001FFC08DFFFFFFFFFBFFC0087FFFFFFFEBF;
defparam dpb_inst_5.INIT_RAM_2D = 256'hFCFFFFFFFFFFFFFFFC27FFFFFFFFFFFFFC08FFFFFFFFFFFFFC1DFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0000000000001F;
defparam dpb_inst_5.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

endmodule //blk_mem_gen_4
